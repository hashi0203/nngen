

module test
(

);

  reg CLK;
  reg RESETN;
  wire irq;
  wire [32-1:0] maxi_awaddr;
  wire [8-1:0] maxi_awlen;
  wire [3-1:0] maxi_awsize;
  wire [2-1:0] maxi_awburst;
  wire [1-1:0] maxi_awlock;
  wire [4-1:0] maxi_awcache;
  wire [3-1:0] maxi_awprot;
  wire [4-1:0] maxi_awqos;
  wire [2-1:0] maxi_awuser;
  wire maxi_awvalid;
  reg maxi_awready;
  wire [32-1:0] maxi_wdata;
  wire [4-1:0] maxi_wstrb;
  wire maxi_wlast;
  wire maxi_wvalid;
  reg maxi_wready;
  reg [2-1:0] maxi_bresp;
  reg maxi_bvalid;
  wire maxi_bready;
  wire [32-1:0] maxi_araddr;
  wire [8-1:0] maxi_arlen;
  wire [3-1:0] maxi_arsize;
  wire [2-1:0] maxi_arburst;
  wire [1-1:0] maxi_arlock;
  wire [4-1:0] maxi_arcache;
  wire [3-1:0] maxi_arprot;
  wire [4-1:0] maxi_arqos;
  wire [2-1:0] maxi_aruser;
  wire maxi_arvalid;
  reg maxi_arready;
  reg [32-1:0] maxi_rdata;
  reg [2-1:0] maxi_rresp;
  reg maxi_rlast;
  reg maxi_rvalid;
  wire maxi_rready;
  reg [32-1:0] saxi_awaddr;
  reg [4-1:0] saxi_awcache;
  reg [3-1:0] saxi_awprot;
  reg saxi_awvalid;
  wire saxi_awready;
  reg [32-1:0] saxi_wdata;
  reg [4-1:0] saxi_wstrb;
  reg saxi_wvalid;
  wire saxi_wready;
  wire [2-1:0] saxi_bresp;
  wire saxi_bvalid;
  reg saxi_bready;
  reg [32-1:0] saxi_araddr;
  reg [4-1:0] saxi_arcache;
  reg [3-1:0] saxi_arprot;
  reg saxi_arvalid;
  wire saxi_arready;
  wire [32-1:0] saxi_rdata;
  wire [2-1:0] saxi_rresp;
  wire saxi_rvalid;
  reg saxi_rready;
  wire RST;
  assign RST = !RESETN;
  wire [32-1:0] memory_awaddr;
  wire [8-1:0] memory_awlen;
  wire [3-1:0] memory_awsize;
  wire [2-1:0] memory_awburst;
  wire [1-1:0] memory_awlock;
  wire [4-1:0] memory_awcache;
  wire [3-1:0] memory_awprot;
  wire [4-1:0] memory_awqos;
  wire [2-1:0] memory_awuser;
  wire memory_awvalid;
  reg memory_awready;
  wire [32-1:0] memory_wdata;
  wire [4-1:0] memory_wstrb;
  wire memory_wlast;
  wire memory_wvalid;
  reg memory_wready;
  wire [2-1:0] memory_bresp;
  reg memory_bvalid;
  wire memory_bready;
  wire [32-1:0] memory_araddr;
  wire [8-1:0] memory_arlen;
  wire [3-1:0] memory_arsize;
  wire [2-1:0] memory_arburst;
  wire [1-1:0] memory_arlock;
  wire [4-1:0] memory_arcache;
  wire [3-1:0] memory_arprot;
  wire [4-1:0] memory_arqos;
  wire [2-1:0] memory_aruser;
  wire memory_arvalid;
  reg memory_arready;
  reg [32-1:0] memory_rdata;
  wire [2-1:0] memory_rresp;
  reg memory_rlast;
  reg memory_rvalid;
  wire memory_rready;
  assign memory_bresp = 0;
  assign memory_rresp = 0;
  reg [32-1:0] _memory_waddr_fsm;
  localparam _memory_waddr_fsm_init = 0;
  reg [32-1:0] _memory_wdata_fsm;
  localparam _memory_wdata_fsm_init = 0;
  reg [32-1:0] _memory_raddr_fsm;
  localparam _memory_raddr_fsm_init = 0;
  reg [32-1:0] _memory_rdata_fsm;
  localparam _memory_rdata_fsm_init = 0;
  wire _memory_wreq_fifo_enq;
  wire [41-1:0] _memory_wreq_fifo_wdata;
  wire _memory_wreq_fifo_full;
  wire _memory_wreq_fifo_almost_full;
  wire _memory_wreq_fifo_deq;
  wire [41-1:0] _memory_wreq_fifo_rdata;
  wire _memory_wreq_fifo_empty;
  wire _memory_wreq_fifo_almost_empty;

  _memory_wreq_fifo
  inst__memory_wreq_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._memory_wreq_fifo_enq(_memory_wreq_fifo_enq),
    ._memory_wreq_fifo_wdata(_memory_wreq_fifo_wdata),
    ._memory_wreq_fifo_full(_memory_wreq_fifo_full),
    ._memory_wreq_fifo_almost_full(_memory_wreq_fifo_almost_full),
    ._memory_wreq_fifo_deq(_memory_wreq_fifo_deq),
    ._memory_wreq_fifo_rdata(_memory_wreq_fifo_rdata),
    ._memory_wreq_fifo_empty(_memory_wreq_fifo_empty),
    ._memory_wreq_fifo_almost_empty(_memory_wreq_fifo_almost_empty)
  );

  reg [4-1:0] count__memory_wreq_fifo;
  wire _memory_rreq_fifo_enq;
  wire [41-1:0] _memory_rreq_fifo_wdata;
  wire _memory_rreq_fifo_full;
  wire _memory_rreq_fifo_almost_full;
  wire _memory_rreq_fifo_deq;
  wire [41-1:0] _memory_rreq_fifo_rdata;
  wire _memory_rreq_fifo_empty;
  wire _memory_rreq_fifo_almost_empty;

  _memory_rreq_fifo
  inst__memory_rreq_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._memory_rreq_fifo_enq(_memory_rreq_fifo_enq),
    ._memory_rreq_fifo_wdata(_memory_rreq_fifo_wdata),
    ._memory_rreq_fifo_full(_memory_rreq_fifo_full),
    ._memory_rreq_fifo_almost_full(_memory_rreq_fifo_almost_full),
    ._memory_rreq_fifo_deq(_memory_rreq_fifo_deq),
    ._memory_rreq_fifo_rdata(_memory_rreq_fifo_rdata),
    ._memory_rreq_fifo_empty(_memory_rreq_fifo_empty),
    ._memory_rreq_fifo_almost_empty(_memory_rreq_fifo_almost_empty)
  );

  reg [4-1:0] count__memory_rreq_fifo;
  reg [8-1:0] _memory_mem [0:2**23-1];

  initial begin
    $readmemh("memimg_test_matrix_conv2d_celu_int32_3x3_stride1.out", _memory_mem);
  end

  reg [33-1:0] _write_count;
  reg [32-1:0] _write_addr;
  reg [33-1:0] _read_count;
  reg [32-1:0] _read_addr;
  reg [33-1:0] _sleep_interval_count;
  reg [33-1:0] _keep_sleep_count;
  wire [32-1:0] pack_write_req_global_addr_0;
  wire [9-1:0] pack_write_req_size_1;
  assign pack_write_req_global_addr_0 = memory_awaddr;
  assign pack_write_req_size_1 = memory_awlen + 1;
  wire [41-1:0] pack_write_req_packed_2;
  assign pack_write_req_packed_2 = { pack_write_req_global_addr_0, pack_write_req_size_1 };
  assign _memory_wreq_fifo_wdata = ((_memory_waddr_fsm == 11) && memory_awvalid && memory_awready)? pack_write_req_packed_2 : 'hx;
  assign _memory_wreq_fifo_enq = ((_memory_waddr_fsm == 11) && memory_awvalid && memory_awready)? (_memory_waddr_fsm == 11) && memory_awvalid && memory_awready && !_memory_wreq_fifo_almost_full : 0;
  localparam _tmp_3 = 1;
  wire [_tmp_3-1:0] _tmp_4;
  assign _tmp_4 = !_memory_wreq_fifo_almost_full;
  reg [_tmp_3-1:0] __tmp_4_1;
  wire [32-1:0] unpack_write_req_global_addr_5;
  wire [9-1:0] unpack_write_req_size_6;
  assign unpack_write_req_global_addr_5 = _memory_wreq_fifo_rdata[40:9];
  assign unpack_write_req_size_6 = _memory_wreq_fifo_rdata[8:0];
  assign _memory_wreq_fifo_deq = ((_memory_wdata_fsm == 0) && !_memory_wreq_fifo_empty && !_memory_wreq_fifo_empty)? 1 : 0;
  wire [32-1:0] pack_read_req_global_addr_7;
  wire [9-1:0] pack_read_req_size_8;
  assign pack_read_req_global_addr_7 = memory_araddr;
  assign pack_read_req_size_8 = memory_arlen + 1;
  wire [41-1:0] pack_read_req_packed_9;
  assign pack_read_req_packed_9 = { pack_read_req_global_addr_7, pack_read_req_size_8 };
  assign _memory_rreq_fifo_wdata = ((_memory_raddr_fsm == 1) && memory_arvalid && memory_arready)? pack_read_req_packed_9 : 'hx;
  assign _memory_rreq_fifo_enq = ((_memory_raddr_fsm == 1) && memory_arvalid && memory_arready)? (_memory_raddr_fsm == 1) && memory_arvalid && memory_arready && !_memory_rreq_fifo_almost_full : 0;
  localparam _tmp_10 = 1;
  wire [_tmp_10-1:0] _tmp_11;
  assign _tmp_11 = !_memory_rreq_fifo_almost_full;
  reg [_tmp_10-1:0] __tmp_11_1;
  wire [32-1:0] unpack_read_req_global_addr_12;
  wire [9-1:0] unpack_read_req_size_13;
  assign unpack_read_req_global_addr_12 = _memory_rreq_fifo_rdata[40:9];
  assign unpack_read_req_size_13 = _memory_rreq_fifo_rdata[8:0];
  assign _memory_rreq_fifo_deq = ((_memory_rdata_fsm == 0) && !_memory_rreq_fifo_empty && !_memory_rreq_fifo_empty)? 1 : 0;
  reg [32-1:0] _d1__memory_rdata_fsm;
  reg __memory_rdata_fsm_cond_11_0_1;
  assign memory_awaddr = maxi_awaddr;
  assign memory_awlen = maxi_awlen;
  assign memory_awsize = maxi_awsize;
  assign memory_awburst = maxi_awburst;
  assign memory_awlock = maxi_awlock;
  assign memory_awcache = maxi_awcache;
  assign memory_awprot = maxi_awprot;
  assign memory_awqos = maxi_awqos;
  assign memory_awuser = maxi_awuser;
  assign memory_awvalid = maxi_awvalid;
  wire _tmp_14;
  assign _tmp_14 = memory_awready;

  always @(*) begin
    maxi_awready = _tmp_14;
  end

  assign memory_wdata = maxi_wdata;
  assign memory_wstrb = maxi_wstrb;
  assign memory_wlast = maxi_wlast;
  assign memory_wvalid = maxi_wvalid;
  wire _tmp_15;
  assign _tmp_15 = memory_wready;

  always @(*) begin
    maxi_wready = _tmp_15;
  end

  wire [2-1:0] _tmp_16;
  assign _tmp_16 = memory_bresp;

  always @(*) begin
    maxi_bresp = _tmp_16;
  end

  wire _tmp_17;
  assign _tmp_17 = memory_bvalid;

  always @(*) begin
    maxi_bvalid = _tmp_17;
  end

  assign memory_bready = maxi_bready;
  assign memory_araddr = maxi_araddr;
  assign memory_arlen = maxi_arlen;
  assign memory_arsize = maxi_arsize;
  assign memory_arburst = maxi_arburst;
  assign memory_arlock = maxi_arlock;
  assign memory_arcache = maxi_arcache;
  assign memory_arprot = maxi_arprot;
  assign memory_arqos = maxi_arqos;
  assign memory_aruser = maxi_aruser;
  assign memory_arvalid = maxi_arvalid;
  wire _tmp_18;
  assign _tmp_18 = memory_arready;

  always @(*) begin
    maxi_arready = _tmp_18;
  end

  wire [32-1:0] _tmp_19;
  assign _tmp_19 = memory_rdata;

  always @(*) begin
    maxi_rdata = _tmp_19;
  end

  wire [2-1:0] _tmp_20;
  assign _tmp_20 = memory_rresp;

  always @(*) begin
    maxi_rresp = _tmp_20;
  end

  wire _tmp_21;
  assign _tmp_21 = memory_rlast;

  always @(*) begin
    maxi_rlast = _tmp_21;
  end

  wire _tmp_22;
  assign _tmp_22 = memory_rvalid;

  always @(*) begin
    maxi_rvalid = _tmp_22;
  end

  assign memory_rready = maxi_rready;
  reg [32-1:0] _saxi_awaddr;
  wire [4-1:0] _saxi_awcache;
  wire [3-1:0] _saxi_awprot;
  reg _saxi_awvalid;
  wire _saxi_awready;
  reg [32-1:0] _saxi_wdata;
  reg [4-1:0] _saxi_wstrb;
  reg _saxi_wvalid;
  wire _saxi_wready;
  wire [2-1:0] _saxi_bresp;
  wire _saxi_bvalid;
  wire _saxi_bready;
  reg [32-1:0] _saxi_araddr;
  wire [4-1:0] _saxi_arcache;
  wire [3-1:0] _saxi_arprot;
  reg _saxi_arvalid;
  wire _saxi_arready;
  wire [32-1:0] _saxi_rdata;
  wire [2-1:0] _saxi_rresp;
  wire _saxi_rvalid;
  wire _saxi_rready;
  assign _saxi_awcache = 3;
  assign _saxi_awprot = 0;
  assign _saxi_bready = 1;
  assign _saxi_arcache = 3;
  assign _saxi_arprot = 0;
  reg [3-1:0] outstanding_wcount_23;
  wire [32-1:0] _tmp_24;
  assign _tmp_24 = _saxi_awaddr;

  always @(*) begin
    saxi_awaddr = _tmp_24;
  end

  wire [4-1:0] _tmp_25;
  assign _tmp_25 = _saxi_awcache;

  always @(*) begin
    saxi_awcache = _tmp_25;
  end

  wire [3-1:0] _tmp_26;
  assign _tmp_26 = _saxi_awprot;

  always @(*) begin
    saxi_awprot = _tmp_26;
  end

  wire _tmp_27;
  assign _tmp_27 = _saxi_awvalid;

  always @(*) begin
    saxi_awvalid = _tmp_27;
  end

  assign _saxi_awready = saxi_awready;
  wire [32-1:0] _tmp_28;
  assign _tmp_28 = _saxi_wdata;

  always @(*) begin
    saxi_wdata = _tmp_28;
  end

  wire [4-1:0] _tmp_29;
  assign _tmp_29 = _saxi_wstrb;

  always @(*) begin
    saxi_wstrb = _tmp_29;
  end

  wire _tmp_30;
  assign _tmp_30 = _saxi_wvalid;

  always @(*) begin
    saxi_wvalid = _tmp_30;
  end

  assign _saxi_wready = saxi_wready;
  assign _saxi_bresp = saxi_bresp;
  assign _saxi_bvalid = saxi_bvalid;
  wire _tmp_31;
  assign _tmp_31 = _saxi_bready;

  always @(*) begin
    saxi_bready = _tmp_31;
  end

  wire [32-1:0] _tmp_32;
  assign _tmp_32 = _saxi_araddr;

  always @(*) begin
    saxi_araddr = _tmp_32;
  end

  wire [4-1:0] _tmp_33;
  assign _tmp_33 = _saxi_arcache;

  always @(*) begin
    saxi_arcache = _tmp_33;
  end

  wire [3-1:0] _tmp_34;
  assign _tmp_34 = _saxi_arprot;

  always @(*) begin
    saxi_arprot = _tmp_34;
  end

  wire _tmp_35;
  assign _tmp_35 = _saxi_arvalid;

  always @(*) begin
    saxi_arvalid = _tmp_35;
  end

  assign _saxi_arready = saxi_arready;
  assign _saxi_rdata = saxi_rdata;
  assign _saxi_rresp = saxi_rresp;
  assign _saxi_rvalid = saxi_rvalid;
  wire _tmp_36;
  assign _tmp_36 = _saxi_rready;

  always @(*) begin
    saxi_rready = _tmp_36;
  end

  reg [32-1:0] time_counter;
  reg [32-1:0] th_ctrl;
  localparam th_ctrl_init = 0;
  reg signed [32-1:0] _th_ctrl_i_0;
  reg __saxi_cond_0_1;
  reg __saxi_cond_1_1;
  reg signed [32-1:0] _th_ctrl_start_time_1;
  reg __saxi_cond_2_1;
  reg __saxi_cond_3_1;
  reg __saxi_cond_4_1;
  reg signed [32-1:0] axim_rdata_37;
  reg __saxi_cond_5_1;
  reg signed [32-1:0] axim_rdata_38;
  assign _saxi_rready = (th_ctrl == 13) || (th_ctrl == 18);
  reg signed [32-1:0] _th_ctrl_end_time_2;
  reg signed [32-1:0] _th_ctrl_ok_3;
  reg signed [32-1:0] _th_ctrl_bat_4;
  reg signed [32-1:0] _th_ctrl_y_5;
  reg signed [32-1:0] _th_ctrl_x_6;
  reg signed [32-1:0] _th_ctrl_ch_7;
  reg signed [32-1:0] rdata_39;
  reg signed [32-1:0] _th_ctrl_orig_8;
  reg signed [32-1:0] rdata_40;
  reg signed [32-1:0] _th_ctrl_check_9;

  matrix_conv2d_celu
  uut
  (
    .CLK(CLK),
    .RESETN(RESETN),
    .irq(irq),
    .maxi_awaddr(maxi_awaddr),
    .maxi_awlen(maxi_awlen),
    .maxi_awsize(maxi_awsize),
    .maxi_awburst(maxi_awburst),
    .maxi_awlock(maxi_awlock),
    .maxi_awcache(maxi_awcache),
    .maxi_awprot(maxi_awprot),
    .maxi_awqos(maxi_awqos),
    .maxi_awuser(maxi_awuser),
    .maxi_awvalid(maxi_awvalid),
    .maxi_awready(maxi_awready),
    .maxi_wdata(maxi_wdata),
    .maxi_wstrb(maxi_wstrb),
    .maxi_wlast(maxi_wlast),
    .maxi_wvalid(maxi_wvalid),
    .maxi_wready(maxi_wready),
    .maxi_bresp(maxi_bresp),
    .maxi_bvalid(maxi_bvalid),
    .maxi_bready(maxi_bready),
    .maxi_araddr(maxi_araddr),
    .maxi_arlen(maxi_arlen),
    .maxi_arsize(maxi_arsize),
    .maxi_arburst(maxi_arburst),
    .maxi_arlock(maxi_arlock),
    .maxi_arcache(maxi_arcache),
    .maxi_arprot(maxi_arprot),
    .maxi_arqos(maxi_arqos),
    .maxi_aruser(maxi_aruser),
    .maxi_arvalid(maxi_arvalid),
    .maxi_arready(maxi_arready),
    .maxi_rdata(maxi_rdata),
    .maxi_rresp(maxi_rresp),
    .maxi_rlast(maxi_rlast),
    .maxi_rvalid(maxi_rvalid),
    .maxi_rready(maxi_rready),
    .saxi_awaddr(saxi_awaddr),
    .saxi_awcache(saxi_awcache),
    .saxi_awprot(saxi_awprot),
    .saxi_awvalid(saxi_awvalid),
    .saxi_awready(saxi_awready),
    .saxi_wdata(saxi_wdata),
    .saxi_wstrb(saxi_wstrb),
    .saxi_wvalid(saxi_wvalid),
    .saxi_wready(saxi_wready),
    .saxi_bresp(saxi_bresp),
    .saxi_bvalid(saxi_bvalid),
    .saxi_bready(saxi_bready),
    .saxi_araddr(saxi_araddr),
    .saxi_arcache(saxi_arcache),
    .saxi_arprot(saxi_arprot),
    .saxi_arvalid(saxi_arvalid),
    .saxi_arready(saxi_arready),
    .saxi_rdata(saxi_rdata),
    .saxi_rresp(saxi_rresp),
    .saxi_rvalid(saxi_rvalid),
    .saxi_rready(saxi_rready)
  );


  initial begin
    CLK = 0;
    forever begin
      #5 CLK = !CLK;
    end
  end


  initial begin
    RESETN = 1;
    memory_awready = 0;
    memory_wready = 0;
    memory_bvalid = 0;
    memory_arready = 0;
    memory_rdata = 0;
    memory_rlast = 0;
    memory_rvalid = 0;
    _memory_waddr_fsm = _memory_waddr_fsm_init;
    _memory_wdata_fsm = _memory_wdata_fsm_init;
    _memory_raddr_fsm = _memory_raddr_fsm_init;
    _memory_rdata_fsm = _memory_rdata_fsm_init;
    count__memory_wreq_fifo = 0;
    count__memory_rreq_fifo = 0;
    _write_count = 0;
    _write_addr = 0;
    _read_count = 0;
    _read_addr = 0;
    _sleep_interval_count = 0;
    _keep_sleep_count = 0;
    __tmp_4_1 = 0;
    __tmp_11_1 = 0;
    _d1__memory_rdata_fsm = _memory_rdata_fsm_init;
    __memory_rdata_fsm_cond_11_0_1 = 0;
    _saxi_awaddr = 0;
    _saxi_awvalid = 0;
    _saxi_wdata = 0;
    _saxi_wstrb = 0;
    _saxi_wvalid = 0;
    _saxi_araddr = 0;
    _saxi_arvalid = 0;
    outstanding_wcount_23 = 0;
    time_counter = 0;
    th_ctrl = th_ctrl_init;
    _th_ctrl_i_0 = 0;
    __saxi_cond_0_1 = 0;
    __saxi_cond_1_1 = 0;
    _th_ctrl_start_time_1 = 0;
    __saxi_cond_2_1 = 0;
    __saxi_cond_3_1 = 0;
    __saxi_cond_4_1 = 0;
    axim_rdata_37 = 0;
    __saxi_cond_5_1 = 0;
    axim_rdata_38 = 0;
    _th_ctrl_end_time_2 = 0;
    _th_ctrl_ok_3 = 0;
    _th_ctrl_bat_4 = 0;
    _th_ctrl_y_5 = 0;
    _th_ctrl_x_6 = 0;
    _th_ctrl_ch_7 = 0;
    rdata_39 = 0;
    _th_ctrl_orig_8 = 0;
    rdata_40 = 0;
    _th_ctrl_check_9 = 0;
    #100;
    RESETN = 0;
    #100;
    RESETN = 1;
    #10000000;
    $finish;
  end


  always @(posedge CLK) begin
    if(RST) begin
      _keep_sleep_count <= 0;
      _sleep_interval_count <= 0;
    end else begin
      if(_sleep_interval_count == 15) begin
        _keep_sleep_count <= _keep_sleep_count + 1;
      end 
      if((_sleep_interval_count == 15) && (_keep_sleep_count == 3)) begin
        _keep_sleep_count <= 0;
      end 
      if(_sleep_interval_count < 15) begin
        _sleep_interval_count <= _sleep_interval_count + 1;
      end 
      if((_keep_sleep_count == 3) && (_sleep_interval_count == 15)) begin
        _sleep_interval_count <= 0;
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[0]) begin
        _memory_mem[_write_addr + 0] <= memory_wdata[7:0];
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[1]) begin
        _memory_mem[_write_addr + 1] <= memory_wdata[15:8];
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[2]) begin
        _memory_mem[_write_addr + 2] <= memory_wdata[23:16];
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[3]) begin
        _memory_mem[_write_addr + 3] <= memory_wdata[31:24];
      end 
    end
  end

  localparam _memory_waddr_fsm_1 = 1;
  localparam _memory_waddr_fsm_2 = 2;
  localparam _memory_waddr_fsm_3 = 3;
  localparam _memory_waddr_fsm_4 = 4;
  localparam _memory_waddr_fsm_5 = 5;
  localparam _memory_waddr_fsm_6 = 6;
  localparam _memory_waddr_fsm_7 = 7;
  localparam _memory_waddr_fsm_8 = 8;
  localparam _memory_waddr_fsm_9 = 9;
  localparam _memory_waddr_fsm_10 = 10;
  localparam _memory_waddr_fsm_11 = 11;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_waddr_fsm <= _memory_waddr_fsm_init;
      memory_awready <= 0;
    end else begin
      case(_memory_waddr_fsm)
        _memory_waddr_fsm_init: begin
          memory_awready <= 0;
          if(memory_awvalid) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_1;
          end 
        end
        _memory_waddr_fsm_1: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_2;
        end
        _memory_waddr_fsm_2: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_3;
        end
        _memory_waddr_fsm_3: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_4;
        end
        _memory_waddr_fsm_4: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_5;
        end
        _memory_waddr_fsm_5: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_6;
        end
        _memory_waddr_fsm_6: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_7;
        end
        _memory_waddr_fsm_7: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_8;
        end
        _memory_waddr_fsm_8: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_9;
        end
        _memory_waddr_fsm_9: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_10;
        end
        _memory_waddr_fsm_10: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_11;
        end
        _memory_waddr_fsm_11: begin
          if(!_memory_wreq_fifo_almost_full) begin
            memory_awready <= 1;
          end 
          if(memory_awvalid && memory_awready) begin
            memory_awready <= 0;
          end 
          if(!memory_awvalid) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_init;
          end 
          if(memory_awvalid && memory_awready) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_wdata_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_wdata_fsm <= _memory_wdata_fsm_init;
      memory_bvalid <= 0;
      _write_addr <= 0;
      _write_count <= 0;
      memory_wready <= 0;
    end else begin
      case(_memory_wdata_fsm)
        _memory_wdata_fsm_init: begin
          memory_bvalid <= 0;
          if(!_memory_wreq_fifo_empty) begin
            _write_addr <= unpack_write_req_global_addr_5;
            _write_count <= unpack_write_req_size_6;
            memory_wready <= 1;
          end 
          if(!_memory_wreq_fifo_empty) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_1;
          end 
        end
        _memory_wdata_fsm_1: begin
          if(memory_wvalid && memory_wready) begin
            _write_addr <= _write_addr + 4;
            _write_count <= _write_count - 1;
          end 
          if(_sleep_interval_count == 15) begin
            memory_wready <= 0;
          end else begin
            memory_wready <= 1;
          end
          if(memory_wvalid && memory_wready && (_write_count == 1)) begin
            memory_wready <= 0;
            memory_bvalid <= 1;
          end 
          if(memory_wvalid && memory_wready && memory_wlast) begin
            memory_wready <= 0;
            memory_bvalid <= 1;
          end 
          if(memory_wvalid && memory_wready && (_write_count == 1)) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_init;
          end 
          if(memory_wvalid && memory_wready && memory_wlast) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_raddr_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_raddr_fsm <= _memory_raddr_fsm_init;
      memory_arready <= 0;
    end else begin
      case(_memory_raddr_fsm)
        _memory_raddr_fsm_init: begin
          memory_arready <= 0;
          if(memory_arvalid) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_1;
          end 
        end
        _memory_raddr_fsm_1: begin
          if(!_memory_rreq_fifo_almost_full) begin
            memory_arready <= 1;
          end 
          if(memory_arvalid && memory_arready) begin
            memory_arready <= 0;
          end 
          if(!memory_arvalid) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_init;
          end 
          if(memory_arvalid && memory_arready) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_rdata_fsm_1 = 1;
  localparam _memory_rdata_fsm_2 = 2;
  localparam _memory_rdata_fsm_3 = 3;
  localparam _memory_rdata_fsm_4 = 4;
  localparam _memory_rdata_fsm_5 = 5;
  localparam _memory_rdata_fsm_6 = 6;
  localparam _memory_rdata_fsm_7 = 7;
  localparam _memory_rdata_fsm_8 = 8;
  localparam _memory_rdata_fsm_9 = 9;
  localparam _memory_rdata_fsm_10 = 10;
  localparam _memory_rdata_fsm_11 = 11;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_rdata_fsm <= _memory_rdata_fsm_init;
      _d1__memory_rdata_fsm <= _memory_rdata_fsm_init;
      _read_addr <= 0;
      _read_count <= 0;
      memory_rdata[7:0] <= (0 >> 0) & { 8{ 1'd1 } };
      memory_rdata[15:8] <= (0 >> 8) & { 8{ 1'd1 } };
      memory_rdata[23:16] <= (0 >> 16) & { 8{ 1'd1 } };
      memory_rdata[31:24] <= (0 >> 24) & { 8{ 1'd1 } };
      memory_rvalid <= 0;
      memory_rlast <= 0;
      __memory_rdata_fsm_cond_11_0_1 <= 0;
      memory_rdata <= 0;
    end else begin
      _d1__memory_rdata_fsm <= _memory_rdata_fsm;
      case(_d1__memory_rdata_fsm)
        _memory_rdata_fsm_11: begin
          if(__memory_rdata_fsm_cond_11_0_1) begin
            memory_rvalid <= 0;
            memory_rlast <= 0;
          end 
        end
      endcase
      case(_memory_rdata_fsm)
        _memory_rdata_fsm_init: begin
          if(!_memory_rreq_fifo_empty) begin
            _read_addr <= unpack_read_req_global_addr_12;
            _read_count <= unpack_read_req_size_13;
          end 
          if(!_memory_rreq_fifo_empty) begin
            _memory_rdata_fsm <= _memory_rdata_fsm_1;
          end 
        end
        _memory_rdata_fsm_1: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_2;
        end
        _memory_rdata_fsm_2: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_3;
        end
        _memory_rdata_fsm_3: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_4;
        end
        _memory_rdata_fsm_4: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_5;
        end
        _memory_rdata_fsm_5: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_6;
        end
        _memory_rdata_fsm_6: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_7;
        end
        _memory_rdata_fsm_7: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_8;
        end
        _memory_rdata_fsm_8: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_9;
        end
        _memory_rdata_fsm_9: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_10;
        end
        _memory_rdata_fsm_10: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_11;
        end
        _memory_rdata_fsm_11: begin
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[7:0] <= _memory_mem[_read_addr + 0];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[15:8] <= _memory_mem[_read_addr + 1];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[23:16] <= _memory_mem[_read_addr + 2];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[31:24] <= _memory_mem[_read_addr + 3];
          end 
          if((_sleep_interval_count < 15) && (_read_count > 0) && memory_rready | !memory_rvalid) begin
            memory_rvalid <= 1;
            _read_addr <= _read_addr + 4;
            _read_count <= _read_count - 1;
          end 
          if((_sleep_interval_count < 15) && (_read_count == 1) && memory_rready | !memory_rvalid) begin
            memory_rlast <= 1;
          end 
          __memory_rdata_fsm_cond_11_0_1 <= 1;
          if(memory_rvalid && !memory_rready) begin
            memory_rvalid <= memory_rvalid;
            memory_rdata <= memory_rdata;
            memory_rlast <= memory_rlast;
          end 
          if(memory_rvalid && memory_rready && (_read_count == 0)) begin
            _memory_rdata_fsm <= _memory_rdata_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__memory_wreq_fifo <= 0;
      __tmp_4_1 <= 0;
    end else begin
      if(_memory_wreq_fifo_enq && !_memory_wreq_fifo_full && (_memory_wreq_fifo_deq && !_memory_wreq_fifo_empty)) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo;
      end else if(_memory_wreq_fifo_enq && !_memory_wreq_fifo_full) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo + 1;
      end else if(_memory_wreq_fifo_deq && !_memory_wreq_fifo_empty) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo - 1;
      end 
      __tmp_4_1 <= _tmp_4;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__memory_rreq_fifo <= 0;
      __tmp_11_1 <= 0;
    end else begin
      if(_memory_rreq_fifo_enq && !_memory_rreq_fifo_full && (_memory_rreq_fifo_deq && !_memory_rreq_fifo_empty)) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo;
      end else if(_memory_rreq_fifo_enq && !_memory_rreq_fifo_full) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo + 1;
      end else if(_memory_rreq_fifo_deq && !_memory_rreq_fifo_empty) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo - 1;
      end 
      __tmp_11_1 <= _tmp_11;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      outstanding_wcount_23 <= 0;
      _saxi_awaddr <= 0;
      _saxi_awvalid <= 0;
      __saxi_cond_0_1 <= 0;
      _saxi_wdata <= 0;
      _saxi_wvalid <= 0;
      _saxi_wstrb <= 0;
      __saxi_cond_1_1 <= 0;
      __saxi_cond_2_1 <= 0;
      __saxi_cond_3_1 <= 0;
      _saxi_araddr <= 0;
      _saxi_arvalid <= 0;
      __saxi_cond_4_1 <= 0;
      __saxi_cond_5_1 <= 0;
    end else begin
      if(__saxi_cond_0_1) begin
        _saxi_awvalid <= 0;
      end 
      if(__saxi_cond_1_1) begin
        _saxi_wvalid <= 0;
      end 
      if(__saxi_cond_2_1) begin
        _saxi_awvalid <= 0;
      end 
      if(__saxi_cond_3_1) begin
        _saxi_wvalid <= 0;
      end 
      if(__saxi_cond_4_1) begin
        _saxi_arvalid <= 0;
      end 
      if(__saxi_cond_5_1) begin
        _saxi_arvalid <= 0;
      end 
      if(_saxi_wvalid && _saxi_wready && !(_saxi_bvalid && _saxi_bready) && (outstanding_wcount_23 < 7)) begin
        outstanding_wcount_23 <= outstanding_wcount_23 + 1;
      end 
      if(!(_saxi_wvalid && _saxi_wready) && (_saxi_bvalid && _saxi_bready) && (outstanding_wcount_23 > 0)) begin
        outstanding_wcount_23 <= outstanding_wcount_23 - 1;
      end 
      if((th_ctrl == 4) && ((outstanding_wcount_23 < 6) && (_saxi_awready || !_saxi_awvalid))) begin
        _saxi_awaddr <= 132;
        _saxi_awvalid <= 1;
      end 
      __saxi_cond_0_1 <= 1;
      if(_saxi_awvalid && !_saxi_awready) begin
        _saxi_awvalid <= _saxi_awvalid;
      end 
      if((th_ctrl == 6) && ((outstanding_wcount_23 < 6) && (_saxi_wready || !_saxi_wvalid))) begin
        _saxi_wdata <= 12544;
        _saxi_wvalid <= 1;
        _saxi_wstrb <= { 4{ 1'd1 } };
      end 
      __saxi_cond_1_1 <= 1;
      if(_saxi_wvalid && !_saxi_wready) begin
        _saxi_wvalid <= _saxi_wvalid;
      end 
      if((th_ctrl == 8) && ((outstanding_wcount_23 < 6) && (_saxi_awready || !_saxi_awvalid))) begin
        _saxi_awaddr <= 16;
        _saxi_awvalid <= 1;
      end 
      __saxi_cond_2_1 <= 1;
      if(_saxi_awvalid && !_saxi_awready) begin
        _saxi_awvalid <= _saxi_awvalid;
      end 
      if((th_ctrl == 10) && ((outstanding_wcount_23 < 6) && (_saxi_wready || !_saxi_wvalid))) begin
        _saxi_wdata <= 1;
        _saxi_wvalid <= 1;
        _saxi_wstrb <= { 4{ 1'd1 } };
      end 
      __saxi_cond_3_1 <= 1;
      if(_saxi_wvalid && !_saxi_wready) begin
        _saxi_wvalid <= _saxi_wvalid;
      end 
      if((th_ctrl == 11) && (_saxi_arready || !_saxi_arvalid)) begin
        _saxi_araddr <= 16;
        _saxi_arvalid <= 1;
      end 
      __saxi_cond_4_1 <= 1;
      if(_saxi_arvalid && !_saxi_arready) begin
        _saxi_arvalid <= _saxi_arvalid;
      end 
      if((th_ctrl == 16) && (_saxi_arready || !_saxi_arvalid)) begin
        _saxi_araddr <= 20;
        _saxi_arvalid <= 1;
      end 
      __saxi_cond_5_1 <= 1;
      if(_saxi_arvalid && !_saxi_arready) begin
        _saxi_arvalid <= _saxi_arvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      time_counter <= 0;
    end else begin
      time_counter <= time_counter + 1;
    end
  end

  localparam th_ctrl_1 = 1;
  localparam th_ctrl_2 = 2;
  localparam th_ctrl_3 = 3;
  localparam th_ctrl_4 = 4;
  localparam th_ctrl_5 = 5;
  localparam th_ctrl_6 = 6;
  localparam th_ctrl_7 = 7;
  localparam th_ctrl_8 = 8;
  localparam th_ctrl_9 = 9;
  localparam th_ctrl_10 = 10;
  localparam th_ctrl_11 = 11;
  localparam th_ctrl_12 = 12;
  localparam th_ctrl_13 = 13;
  localparam th_ctrl_14 = 14;
  localparam th_ctrl_15 = 15;
  localparam th_ctrl_16 = 16;
  localparam th_ctrl_17 = 17;
  localparam th_ctrl_18 = 18;
  localparam th_ctrl_19 = 19;
  localparam th_ctrl_20 = 20;
  localparam th_ctrl_21 = 21;
  localparam th_ctrl_22 = 22;
  localparam th_ctrl_23 = 23;
  localparam th_ctrl_24 = 24;
  localparam th_ctrl_25 = 25;
  localparam th_ctrl_26 = 26;
  localparam th_ctrl_27 = 27;
  localparam th_ctrl_28 = 28;
  localparam th_ctrl_29 = 29;
  localparam th_ctrl_30 = 30;
  localparam th_ctrl_31 = 31;
  localparam th_ctrl_32 = 32;
  localparam th_ctrl_33 = 33;
  localparam th_ctrl_34 = 34;
  localparam th_ctrl_35 = 35;
  localparam th_ctrl_36 = 36;
  localparam th_ctrl_37 = 37;
  localparam th_ctrl_38 = 38;
  localparam th_ctrl_39 = 39;
  localparam th_ctrl_40 = 40;
  localparam th_ctrl_41 = 41;
  localparam th_ctrl_42 = 42;
  localparam th_ctrl_43 = 43;
  localparam th_ctrl_44 = 44;
  localparam th_ctrl_45 = 45;
  localparam th_ctrl_46 = 46;
  localparam th_ctrl_47 = 47;
  localparam th_ctrl_48 = 48;

  always @(posedge CLK) begin
    if(RST) begin
      th_ctrl <= th_ctrl_init;
      _th_ctrl_i_0 <= 0;
      _th_ctrl_start_time_1 <= 0;
      axim_rdata_37 <= 0;
      axim_rdata_38 <= 0;
      _th_ctrl_end_time_2 <= 0;
      _th_ctrl_ok_3 <= 0;
      _th_ctrl_bat_4 <= 0;
      _th_ctrl_y_5 <= 0;
      _th_ctrl_x_6 <= 0;
      _th_ctrl_ch_7 <= 0;
      rdata_39 <= 0;
      _th_ctrl_orig_8 <= 0;
      rdata_40 <= 0;
      _th_ctrl_check_9 <= 0;
    end else begin
      case(th_ctrl)
        th_ctrl_init: begin
          th_ctrl <= th_ctrl_1;
        end
        th_ctrl_1: begin
          _th_ctrl_i_0 <= 0;
          th_ctrl <= th_ctrl_2;
        end
        th_ctrl_2: begin
          if(_th_ctrl_i_0 < 100) begin
            th_ctrl <= th_ctrl_3;
          end else begin
            th_ctrl <= th_ctrl_4;
          end
        end
        th_ctrl_3: begin
          _th_ctrl_i_0 <= _th_ctrl_i_0 + 1;
          th_ctrl <= th_ctrl_2;
        end
        th_ctrl_4: begin
          if((outstanding_wcount_23 < 6) && (_saxi_awready || !_saxi_awvalid)) begin
            th_ctrl <= th_ctrl_5;
          end 
        end
        th_ctrl_5: begin
          th_ctrl <= th_ctrl_6;
        end
        th_ctrl_6: begin
          if(_saxi_wready || !_saxi_wvalid) begin
            th_ctrl <= th_ctrl_7;
          end 
        end
        th_ctrl_7: begin
          _th_ctrl_start_time_1 <= time_counter;
          th_ctrl <= th_ctrl_8;
        end
        th_ctrl_8: begin
          if((outstanding_wcount_23 < 6) && (_saxi_awready || !_saxi_awvalid)) begin
            th_ctrl <= th_ctrl_9;
          end 
        end
        th_ctrl_9: begin
          th_ctrl <= th_ctrl_10;
        end
        th_ctrl_10: begin
          if(_saxi_wready || !_saxi_wvalid) begin
            th_ctrl <= th_ctrl_11;
          end 
        end
        th_ctrl_11: begin
          if(_saxi_arready || !_saxi_arvalid) begin
            th_ctrl <= th_ctrl_12;
          end 
        end
        th_ctrl_12: begin
          th_ctrl <= th_ctrl_13;
        end
        th_ctrl_13: begin
          if(_saxi_rvalid) begin
            axim_rdata_37 <= _saxi_rdata;
          end 
          if(_saxi_rvalid) begin
            th_ctrl <= th_ctrl_14;
          end 
        end
        th_ctrl_14: begin
          if(axim_rdata_37 != 0) begin
            th_ctrl <= th_ctrl_11;
          end 
          if(axim_rdata_37 == 0) begin
            th_ctrl <= th_ctrl_15;
          end 
        end
        th_ctrl_15: begin
          $display("# start");
          th_ctrl <= th_ctrl_16;
        end
        th_ctrl_16: begin
          if(_saxi_arready || !_saxi_arvalid) begin
            th_ctrl <= th_ctrl_17;
          end 
        end
        th_ctrl_17: begin
          th_ctrl <= th_ctrl_18;
        end
        th_ctrl_18: begin
          if(_saxi_rvalid) begin
            axim_rdata_38 <= _saxi_rdata;
          end 
          if(_saxi_rvalid) begin
            th_ctrl <= th_ctrl_19;
          end 
        end
        th_ctrl_19: begin
          if(axim_rdata_38 != 0) begin
            th_ctrl <= th_ctrl_16;
          end 
          if(axim_rdata_38 == 0) begin
            th_ctrl <= th_ctrl_20;
          end 
        end
        th_ctrl_20: begin
          _th_ctrl_end_time_2 <= time_counter;
          th_ctrl <= th_ctrl_21;
        end
        th_ctrl_21: begin
          $display("# end");
          th_ctrl <= th_ctrl_22;
        end
        th_ctrl_22: begin
          $display("# execution cycles: %d", (_th_ctrl_end_time_2 - _th_ctrl_start_time_1));
          th_ctrl <= th_ctrl_23;
        end
        th_ctrl_23: begin
          _th_ctrl_ok_3 <= 1;
          th_ctrl <= th_ctrl_24;
        end
        th_ctrl_24: begin
          _th_ctrl_bat_4 <= 0;
          th_ctrl <= th_ctrl_25;
        end
        th_ctrl_25: begin
          if(_th_ctrl_bat_4 < 1) begin
            th_ctrl <= th_ctrl_26;
          end else begin
            th_ctrl <= th_ctrl_43;
          end
        end
        th_ctrl_26: begin
          _th_ctrl_y_5 <= 0;
          th_ctrl <= th_ctrl_27;
        end
        th_ctrl_27: begin
          if(_th_ctrl_y_5 < 7) begin
            th_ctrl <= th_ctrl_28;
          end else begin
            th_ctrl <= th_ctrl_42;
          end
        end
        th_ctrl_28: begin
          _th_ctrl_x_6 <= 0;
          th_ctrl <= th_ctrl_29;
        end
        th_ctrl_29: begin
          if(_th_ctrl_x_6 < 7) begin
            th_ctrl <= th_ctrl_30;
          end else begin
            th_ctrl <= th_ctrl_41;
          end
        end
        th_ctrl_30: begin
          _th_ctrl_ch_7 <= 0;
          th_ctrl <= th_ctrl_31;
        end
        th_ctrl_31: begin
          if(_th_ctrl_ch_7 < 7) begin
            th_ctrl <= th_ctrl_32;
          end else begin
            th_ctrl <= th_ctrl_40;
          end
        end
        th_ctrl_32: begin
          if(th_ctrl == 32) begin
            rdata_39 <= { _memory_mem[0 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 3], _memory_mem[0 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 2], _memory_mem[0 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 1], _memory_mem[0 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 0] } >> (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 % 8;
          end 
          th_ctrl <= th_ctrl_33;
        end
        th_ctrl_33: begin
          _th_ctrl_orig_8 <= rdata_39;
          th_ctrl <= th_ctrl_34;
        end
        th_ctrl_34: begin
          if(th_ctrl == 34) begin
            rdata_40 <= { _memory_mem[8448 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 3], _memory_mem[8448 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 2], _memory_mem[8448 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 1], _memory_mem[8448 + (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 / 8 + 0] } >> (_th_ctrl_bat_4 * 7 * 7 * 7 + _th_ctrl_y_5 * 7 * 7 + _th_ctrl_x_6 * 7 + _th_ctrl_ch_7) * 32 % 8;
          end 
          th_ctrl <= th_ctrl_35;
        end
        th_ctrl_35: begin
          _th_ctrl_check_9 <= rdata_40;
          th_ctrl <= th_ctrl_36;
        end
        th_ctrl_36: begin
          if(_th_ctrl_orig_8 !== _th_ctrl_check_9) begin
            th_ctrl <= th_ctrl_37;
          end else begin
            th_ctrl <= th_ctrl_39;
          end
        end
        th_ctrl_37: begin
          $display("NG ( %d %d %d %d ) orig:  %d  check:  %d", _th_ctrl_bat_4, _th_ctrl_y_5, _th_ctrl_x_6, _th_ctrl_ch_7, _th_ctrl_orig_8, _th_ctrl_check_9);
          th_ctrl <= th_ctrl_38;
        end
        th_ctrl_38: begin
          _th_ctrl_ok_3 <= 0;
          th_ctrl <= th_ctrl_39;
        end
        th_ctrl_39: begin
          _th_ctrl_ch_7 <= _th_ctrl_ch_7 + 1;
          th_ctrl <= th_ctrl_31;
        end
        th_ctrl_40: begin
          _th_ctrl_x_6 <= _th_ctrl_x_6 + 1;
          th_ctrl <= th_ctrl_29;
        end
        th_ctrl_41: begin
          _th_ctrl_y_5 <= _th_ctrl_y_5 + 1;
          th_ctrl <= th_ctrl_27;
        end
        th_ctrl_42: begin
          _th_ctrl_bat_4 <= _th_ctrl_bat_4 + 1;
          th_ctrl <= th_ctrl_25;
        end
        th_ctrl_43: begin
          if(_th_ctrl_ok_3) begin
            th_ctrl <= th_ctrl_44;
          end else begin
            th_ctrl <= th_ctrl_46;
          end
        end
        th_ctrl_44: begin
          $display("# verify: PASSED");
          th_ctrl <= th_ctrl_45;
        end
        th_ctrl_45: begin
          th_ctrl <= th_ctrl_47;
        end
        th_ctrl_46: begin
          $display("# verify: FAILED");
          th_ctrl <= th_ctrl_47;
        end
        th_ctrl_47: begin
          $finish;
          th_ctrl <= th_ctrl_48;
        end
      endcase
    end
  end


endmodule



module _memory_wreq_fifo
(
  input CLK,
  input RST,
  input _memory_wreq_fifo_enq,
  input [41-1:0] _memory_wreq_fifo_wdata,
  output _memory_wreq_fifo_full,
  output _memory_wreq_fifo_almost_full,
  input _memory_wreq_fifo_deq,
  output [41-1:0] _memory_wreq_fifo_rdata,
  output _memory_wreq_fifo_empty,
  output _memory_wreq_fifo_almost_empty
);

  reg [41-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [41-1:0] rdata;
  assign _memory_wreq_fifo_full = is_full;
  assign _memory_wreq_fifo_almost_full = is_almost_full || is_full;
  assign _memory_wreq_fifo_empty = is_empty;
  assign _memory_wreq_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _memory_wreq_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_memory_wreq_fifo_enq && !is_full) begin
        mem[head] <= _memory_wreq_fifo_wdata;
        head <= head + 1;
      end 
      if(_memory_wreq_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _memory_rreq_fifo
(
  input CLK,
  input RST,
  input _memory_rreq_fifo_enq,
  input [41-1:0] _memory_rreq_fifo_wdata,
  output _memory_rreq_fifo_full,
  output _memory_rreq_fifo_almost_full,
  input _memory_rreq_fifo_deq,
  output [41-1:0] _memory_rreq_fifo_rdata,
  output _memory_rreq_fifo_empty,
  output _memory_rreq_fifo_almost_empty
);

  reg [41-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [41-1:0] rdata;
  assign _memory_rreq_fifo_full = is_full;
  assign _memory_rreq_fifo_almost_full = is_almost_full || is_full;
  assign _memory_rreq_fifo_empty = is_empty;
  assign _memory_rreq_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _memory_rreq_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_memory_rreq_fifo_enq && !is_full) begin
        mem[head] <= _memory_rreq_fifo_wdata;
        head <= head + 1;
      end 
      if(_memory_rreq_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module matrix_conv2d_celu
(
  input CLK,
  input RESETN,
  output reg irq,
  output reg [32-1:0] maxi_awaddr,
  output reg [8-1:0] maxi_awlen,
  output [3-1:0] maxi_awsize,
  output [2-1:0] maxi_awburst,
  output [1-1:0] maxi_awlock,
  output [4-1:0] maxi_awcache,
  output [3-1:0] maxi_awprot,
  output [4-1:0] maxi_awqos,
  output [2-1:0] maxi_awuser,
  output reg maxi_awvalid,
  input maxi_awready,
  output reg [32-1:0] maxi_wdata,
  output reg [4-1:0] maxi_wstrb,
  output reg maxi_wlast,
  output reg maxi_wvalid,
  input maxi_wready,
  input [2-1:0] maxi_bresp,
  input maxi_bvalid,
  output maxi_bready,
  output reg [32-1:0] maxi_araddr,
  output reg [8-1:0] maxi_arlen,
  output [3-1:0] maxi_arsize,
  output [2-1:0] maxi_arburst,
  output [1-1:0] maxi_arlock,
  output [4-1:0] maxi_arcache,
  output [3-1:0] maxi_arprot,
  output [4-1:0] maxi_arqos,
  output [2-1:0] maxi_aruser,
  output reg maxi_arvalid,
  input maxi_arready,
  input [32-1:0] maxi_rdata,
  input [2-1:0] maxi_rresp,
  input maxi_rlast,
  input maxi_rvalid,
  output maxi_rready,
  input [32-1:0] saxi_awaddr,
  input [4-1:0] saxi_awcache,
  input [3-1:0] saxi_awprot,
  input saxi_awvalid,
  output saxi_awready,
  input [32-1:0] saxi_wdata,
  input [4-1:0] saxi_wstrb,
  input saxi_wvalid,
  output saxi_wready,
  output [2-1:0] saxi_bresp,
  output reg saxi_bvalid,
  input saxi_bready,
  input [32-1:0] saxi_araddr,
  input [4-1:0] saxi_arcache,
  input [3-1:0] saxi_arprot,
  input saxi_arvalid,
  output saxi_arready,
  output reg [32-1:0] saxi_rdata,
  output [2-1:0] saxi_rresp,
  output reg saxi_rvalid,
  input saxi_rready
);

  wire RESETN_inv;
  assign RESETN_inv = !RESETN;
  wire RESETN_inv_buf;
  reg _RESETN_inv_1;
  reg _RESETN_inv_2;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign maxi_awsize = 2;
  assign maxi_awburst = 1;
  assign maxi_awlock = 0;
  assign maxi_awcache = 3;
  assign maxi_awprot = 0;
  assign maxi_awqos = 0;
  assign maxi_awuser = 0;
  assign maxi_bready = 1;
  assign maxi_arsize = 2;
  assign maxi_arburst = 1;
  assign maxi_arlock = 0;
  assign maxi_arcache = 3;
  assign maxi_arprot = 0;
  assign maxi_arqos = 0;
  assign maxi_aruser = 0;
  reg [3-1:0] outstanding_wcount_0;
  reg _maxi_read_start;
  reg [8-1:0] _maxi_read_op_sel;
  reg [32-1:0] _maxi_read_global_addr;
  reg [33-1:0] _maxi_read_global_size;
  reg [32-1:0] _maxi_read_local_addr;
  reg [32-1:0] _maxi_read_local_stride;
  reg [33-1:0] _maxi_read_local_size;
  reg [32-1:0] _maxi_read_local_blocksize;
  wire _maxi_read_req_fifo_enq;
  wire [137-1:0] _maxi_read_req_fifo_wdata;
  wire _maxi_read_req_fifo_full;
  wire _maxi_read_req_fifo_almost_full;
  wire _maxi_read_req_fifo_deq;
  wire [137-1:0] _maxi_read_req_fifo_rdata;
  wire _maxi_read_req_fifo_empty;
  wire _maxi_read_req_fifo_almost_empty;

  _maxi_read_req_fifo
  inst__maxi_read_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_read_req_fifo_enq(_maxi_read_req_fifo_enq),
    ._maxi_read_req_fifo_wdata(_maxi_read_req_fifo_wdata),
    ._maxi_read_req_fifo_full(_maxi_read_req_fifo_full),
    ._maxi_read_req_fifo_almost_full(_maxi_read_req_fifo_almost_full),
    ._maxi_read_req_fifo_deq(_maxi_read_req_fifo_deq),
    ._maxi_read_req_fifo_rdata(_maxi_read_req_fifo_rdata),
    ._maxi_read_req_fifo_empty(_maxi_read_req_fifo_empty),
    ._maxi_read_req_fifo_almost_empty(_maxi_read_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_read_req_fifo;
  wire [8-1:0] _maxi_read_op_sel_fifo;
  wire [32-1:0] _maxi_read_local_addr_fifo;
  wire [32-1:0] _maxi_read_local_stride_fifo;
  wire [33-1:0] _maxi_read_local_size_fifo;
  wire [32-1:0] _maxi_read_local_blocksize_fifo;
  wire [8-1:0] unpack_read_req_op_sel_1;
  wire [32-1:0] unpack_read_req_local_addr_2;
  wire [32-1:0] unpack_read_req_local_stride_3;
  wire [33-1:0] unpack_read_req_local_size_4;
  wire [32-1:0] unpack_read_req_local_blocksize_5;
  assign unpack_read_req_op_sel_1 = _maxi_read_req_fifo_rdata[136:129];
  assign unpack_read_req_local_addr_2 = _maxi_read_req_fifo_rdata[128:97];
  assign unpack_read_req_local_stride_3 = _maxi_read_req_fifo_rdata[96:65];
  assign unpack_read_req_local_size_4 = _maxi_read_req_fifo_rdata[64:32];
  assign unpack_read_req_local_blocksize_5 = _maxi_read_req_fifo_rdata[31:0];
  assign _maxi_read_op_sel_fifo = unpack_read_req_op_sel_1;
  assign _maxi_read_local_addr_fifo = unpack_read_req_local_addr_2;
  assign _maxi_read_local_stride_fifo = unpack_read_req_local_stride_3;
  assign _maxi_read_local_size_fifo = unpack_read_req_local_size_4;
  assign _maxi_read_local_blocksize_fifo = unpack_read_req_local_blocksize_5;
  reg [8-1:0] _maxi_read_op_sel_buf;
  reg [32-1:0] _maxi_read_local_addr_buf;
  reg [32-1:0] _maxi_read_local_stride_buf;
  reg [33-1:0] _maxi_read_local_size_buf;
  reg [32-1:0] _maxi_read_local_blocksize_buf;
  reg _maxi_read_req_idle;
  reg _maxi_read_data_idle;
  wire _maxi_read_idle;
  assign _maxi_read_idle = !_maxi_read_start && _maxi_read_req_idle && _maxi_read_req_fifo_empty && _maxi_read_data_idle;
  reg _maxi_write_start;
  reg [8-1:0] _maxi_write_op_sel;
  reg [32-1:0] _maxi_write_global_addr;
  reg [33-1:0] _maxi_write_global_size;
  reg [32-1:0] _maxi_write_local_addr;
  reg [32-1:0] _maxi_write_local_stride;
  reg [33-1:0] _maxi_write_local_size;
  reg [32-1:0] _maxi_write_local_blocksize;
  wire _maxi_write_req_fifo_enq;
  wire [137-1:0] _maxi_write_req_fifo_wdata;
  wire _maxi_write_req_fifo_full;
  wire _maxi_write_req_fifo_almost_full;
  wire _maxi_write_req_fifo_deq;
  wire [137-1:0] _maxi_write_req_fifo_rdata;
  wire _maxi_write_req_fifo_empty;
  wire _maxi_write_req_fifo_almost_empty;

  _maxi_write_req_fifo
  inst__maxi_write_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_write_req_fifo_enq(_maxi_write_req_fifo_enq),
    ._maxi_write_req_fifo_wdata(_maxi_write_req_fifo_wdata),
    ._maxi_write_req_fifo_full(_maxi_write_req_fifo_full),
    ._maxi_write_req_fifo_almost_full(_maxi_write_req_fifo_almost_full),
    ._maxi_write_req_fifo_deq(_maxi_write_req_fifo_deq),
    ._maxi_write_req_fifo_rdata(_maxi_write_req_fifo_rdata),
    ._maxi_write_req_fifo_empty(_maxi_write_req_fifo_empty),
    ._maxi_write_req_fifo_almost_empty(_maxi_write_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_write_req_fifo;
  wire [8-1:0] _maxi_write_op_sel_fifo;
  wire [32-1:0] _maxi_write_local_addr_fifo;
  wire [32-1:0] _maxi_write_local_stride_fifo;
  wire [33-1:0] _maxi_write_size_fifo;
  wire [32-1:0] _maxi_write_local_blocksize_fifo;
  wire [8-1:0] unpack_write_req_op_sel_6;
  wire [32-1:0] unpack_write_req_local_addr_7;
  wire [32-1:0] unpack_write_req_local_stride_8;
  wire [33-1:0] unpack_write_req_size_9;
  wire [32-1:0] unpack_write_req_local_blocksize_10;
  assign unpack_write_req_op_sel_6 = _maxi_write_req_fifo_rdata[136:129];
  assign unpack_write_req_local_addr_7 = _maxi_write_req_fifo_rdata[128:97];
  assign unpack_write_req_local_stride_8 = _maxi_write_req_fifo_rdata[96:65];
  assign unpack_write_req_size_9 = _maxi_write_req_fifo_rdata[64:32];
  assign unpack_write_req_local_blocksize_10 = _maxi_write_req_fifo_rdata[31:0];
  assign _maxi_write_op_sel_fifo = unpack_write_req_op_sel_6;
  assign _maxi_write_local_addr_fifo = unpack_write_req_local_addr_7;
  assign _maxi_write_local_stride_fifo = unpack_write_req_local_stride_8;
  assign _maxi_write_size_fifo = unpack_write_req_size_9;
  assign _maxi_write_local_blocksize_fifo = unpack_write_req_local_blocksize_10;
  reg [8-1:0] _maxi_write_op_sel_buf;
  reg [32-1:0] _maxi_write_local_addr_buf;
  reg [32-1:0] _maxi_write_local_stride_buf;
  reg [33-1:0] _maxi_write_size_buf;
  reg [32-1:0] _maxi_write_local_blocksize_buf;
  reg _maxi_write_req_idle;
  reg _maxi_write_data_idle;
  wire _maxi_write_idle;
  assign _maxi_write_idle = !_maxi_write_start && _maxi_write_req_idle && _maxi_write_req_fifo_empty && _maxi_write_data_idle;
  reg [32-1:0] _maxi_global_base_addr;
  assign saxi_bresp = 0;
  assign saxi_rresp = 0;
  reg signed [32-1:0] _saxi_register_0;
  reg signed [32-1:0] _saxi_register_1;
  reg signed [32-1:0] _saxi_register_2;
  reg signed [32-1:0] _saxi_register_3;
  reg signed [32-1:0] _saxi_register_4;
  reg signed [32-1:0] _saxi_register_5;
  reg signed [32-1:0] _saxi_register_6;
  reg signed [32-1:0] _saxi_register_7;
  reg signed [32-1:0] _saxi_register_8;
  reg signed [32-1:0] _saxi_register_9;
  reg signed [32-1:0] _saxi_register_10;
  reg signed [32-1:0] _saxi_register_11;
  reg signed [32-1:0] _saxi_register_12;
  reg signed [32-1:0] _saxi_register_13;
  reg signed [32-1:0] _saxi_register_14;
  reg signed [32-1:0] _saxi_register_15;
  reg signed [32-1:0] _saxi_register_16;
  reg signed [32-1:0] _saxi_register_17;
  reg signed [32-1:0] _saxi_register_18;
  reg signed [32-1:0] _saxi_register_19;
  reg signed [32-1:0] _saxi_register_20;
  reg signed [32-1:0] _saxi_register_21;
  reg signed [32-1:0] _saxi_register_22;
  reg signed [32-1:0] _saxi_register_23;
  reg signed [32-1:0] _saxi_register_24;
  reg signed [32-1:0] _saxi_register_25;
  reg signed [32-1:0] _saxi_register_26;
  reg signed [32-1:0] _saxi_register_27;
  reg signed [32-1:0] _saxi_register_28;
  reg signed [32-1:0] _saxi_register_29;
  reg signed [32-1:0] _saxi_register_30;
  reg signed [32-1:0] _saxi_register_31;
  reg signed [32-1:0] _saxi_register_32;
  reg signed [32-1:0] _saxi_register_33;
  reg signed [32-1:0] _saxi_register_34;
  reg signed [32-1:0] _saxi_register_35;
  reg signed [32-1:0] _saxi_register_36;
  reg _saxi_flag_0;
  reg _saxi_flag_1;
  reg _saxi_flag_2;
  reg _saxi_flag_3;
  reg _saxi_flag_4;
  reg _saxi_flag_5;
  reg _saxi_flag_6;
  reg _saxi_flag_7;
  reg _saxi_flag_8;
  reg _saxi_flag_9;
  reg _saxi_flag_10;
  reg _saxi_flag_11;
  reg _saxi_flag_12;
  reg _saxi_flag_13;
  reg _saxi_flag_14;
  reg _saxi_flag_15;
  reg _saxi_flag_16;
  reg _saxi_flag_17;
  reg _saxi_flag_18;
  reg _saxi_flag_19;
  reg _saxi_flag_20;
  reg _saxi_flag_21;
  reg _saxi_flag_22;
  reg _saxi_flag_23;
  reg _saxi_flag_24;
  reg _saxi_flag_25;
  reg _saxi_flag_26;
  reg _saxi_flag_27;
  reg _saxi_flag_28;
  reg _saxi_flag_29;
  reg _saxi_flag_30;
  reg _saxi_flag_31;
  reg _saxi_flag_32;
  reg _saxi_flag_33;
  reg _saxi_flag_34;
  reg _saxi_flag_35;
  reg _saxi_flag_36;
  reg signed [32-1:0] _saxi_resetval_0;
  reg signed [32-1:0] _saxi_resetval_1;
  reg signed [32-1:0] _saxi_resetval_2;
  reg signed [32-1:0] _saxi_resetval_3;
  reg signed [32-1:0] _saxi_resetval_4;
  reg signed [32-1:0] _saxi_resetval_5;
  reg signed [32-1:0] _saxi_resetval_6;
  reg signed [32-1:0] _saxi_resetval_7;
  reg signed [32-1:0] _saxi_resetval_8;
  reg signed [32-1:0] _saxi_resetval_9;
  reg signed [32-1:0] _saxi_resetval_10;
  reg signed [32-1:0] _saxi_resetval_11;
  reg signed [32-1:0] _saxi_resetval_12;
  reg signed [32-1:0] _saxi_resetval_13;
  reg signed [32-1:0] _saxi_resetval_14;
  reg signed [32-1:0] _saxi_resetval_15;
  reg signed [32-1:0] _saxi_resetval_16;
  reg signed [32-1:0] _saxi_resetval_17;
  reg signed [32-1:0] _saxi_resetval_18;
  reg signed [32-1:0] _saxi_resetval_19;
  reg signed [32-1:0] _saxi_resetval_20;
  reg signed [32-1:0] _saxi_resetval_21;
  reg signed [32-1:0] _saxi_resetval_22;
  reg signed [32-1:0] _saxi_resetval_23;
  reg signed [32-1:0] _saxi_resetval_24;
  reg signed [32-1:0] _saxi_resetval_25;
  reg signed [32-1:0] _saxi_resetval_26;
  reg signed [32-1:0] _saxi_resetval_27;
  reg signed [32-1:0] _saxi_resetval_28;
  reg signed [32-1:0] _saxi_resetval_29;
  reg signed [32-1:0] _saxi_resetval_30;
  reg signed [32-1:0] _saxi_resetval_31;
  reg signed [32-1:0] _saxi_resetval_32;
  reg signed [32-1:0] _saxi_resetval_33;
  reg signed [32-1:0] _saxi_resetval_34;
  reg signed [32-1:0] _saxi_resetval_35;
  reg signed [32-1:0] _saxi_resetval_36;
  localparam _saxi_maskwidth = 6;
  localparam _saxi_mask = { _saxi_maskwidth{ 1'd1 } };
  localparam _saxi_shift = 2;
  reg [32-1:0] _saxi_register_fsm;
  localparam _saxi_register_fsm_init = 0;
  reg [32-1:0] addr_11;
  reg writevalid_12;
  reg readvalid_13;
  reg prev_awvalid_14;
  reg prev_arvalid_15;
  assign saxi_awready = (_saxi_register_fsm == 0) && (!writevalid_12 && !readvalid_13 && !saxi_bvalid && prev_awvalid_14);
  assign saxi_arready = (_saxi_register_fsm == 0) && (!readvalid_13 && !writevalid_12 && prev_arvalid_15 && !prev_awvalid_14);
  reg [_saxi_maskwidth-1:0] axis_maskaddr_16;
  wire signed [32-1:0] axislite_rdata_17;
  assign axislite_rdata_17 = (axis_maskaddr_16 == 0)? _saxi_register_0 : 
                             (axis_maskaddr_16 == 1)? _saxi_register_1 : 
                             (axis_maskaddr_16 == 2)? _saxi_register_2 : 
                             (axis_maskaddr_16 == 3)? _saxi_register_3 : 
                             (axis_maskaddr_16 == 4)? _saxi_register_4 : 
                             (axis_maskaddr_16 == 5)? _saxi_register_5 : 
                             (axis_maskaddr_16 == 6)? _saxi_register_6 : 
                             (axis_maskaddr_16 == 7)? _saxi_register_7 : 
                             (axis_maskaddr_16 == 8)? _saxi_register_8 : 
                             (axis_maskaddr_16 == 9)? _saxi_register_9 : 
                             (axis_maskaddr_16 == 10)? _saxi_register_10 : 
                             (axis_maskaddr_16 == 11)? _saxi_register_11 : 
                             (axis_maskaddr_16 == 12)? _saxi_register_12 : 
                             (axis_maskaddr_16 == 13)? _saxi_register_13 : 
                             (axis_maskaddr_16 == 14)? _saxi_register_14 : 
                             (axis_maskaddr_16 == 15)? _saxi_register_15 : 
                             (axis_maskaddr_16 == 16)? _saxi_register_16 : 
                             (axis_maskaddr_16 == 17)? _saxi_register_17 : 
                             (axis_maskaddr_16 == 18)? _saxi_register_18 : 
                             (axis_maskaddr_16 == 19)? _saxi_register_19 : 
                             (axis_maskaddr_16 == 20)? _saxi_register_20 : 
                             (axis_maskaddr_16 == 21)? _saxi_register_21 : 
                             (axis_maskaddr_16 == 22)? _saxi_register_22 : 
                             (axis_maskaddr_16 == 23)? _saxi_register_23 : 
                             (axis_maskaddr_16 == 24)? _saxi_register_24 : 
                             (axis_maskaddr_16 == 25)? _saxi_register_25 : 
                             (axis_maskaddr_16 == 26)? _saxi_register_26 : 
                             (axis_maskaddr_16 == 27)? _saxi_register_27 : 
                             (axis_maskaddr_16 == 28)? _saxi_register_28 : 
                             (axis_maskaddr_16 == 29)? _saxi_register_29 : 
                             (axis_maskaddr_16 == 30)? _saxi_register_30 : 
                             (axis_maskaddr_16 == 31)? _saxi_register_31 : 
                             (axis_maskaddr_16 == 32)? _saxi_register_32 : 
                             (axis_maskaddr_16 == 33)? _saxi_register_33 : 
                             (axis_maskaddr_16 == 34)? _saxi_register_34 : 
                             (axis_maskaddr_16 == 35)? _saxi_register_35 : 
                             (axis_maskaddr_16 == 36)? _saxi_register_36 : 'hx;
  wire axislite_flag_18;
  assign axislite_flag_18 = (axis_maskaddr_16 == 0)? _saxi_flag_0 : 
                            (axis_maskaddr_16 == 1)? _saxi_flag_1 : 
                            (axis_maskaddr_16 == 2)? _saxi_flag_2 : 
                            (axis_maskaddr_16 == 3)? _saxi_flag_3 : 
                            (axis_maskaddr_16 == 4)? _saxi_flag_4 : 
                            (axis_maskaddr_16 == 5)? _saxi_flag_5 : 
                            (axis_maskaddr_16 == 6)? _saxi_flag_6 : 
                            (axis_maskaddr_16 == 7)? _saxi_flag_7 : 
                            (axis_maskaddr_16 == 8)? _saxi_flag_8 : 
                            (axis_maskaddr_16 == 9)? _saxi_flag_9 : 
                            (axis_maskaddr_16 == 10)? _saxi_flag_10 : 
                            (axis_maskaddr_16 == 11)? _saxi_flag_11 : 
                            (axis_maskaddr_16 == 12)? _saxi_flag_12 : 
                            (axis_maskaddr_16 == 13)? _saxi_flag_13 : 
                            (axis_maskaddr_16 == 14)? _saxi_flag_14 : 
                            (axis_maskaddr_16 == 15)? _saxi_flag_15 : 
                            (axis_maskaddr_16 == 16)? _saxi_flag_16 : 
                            (axis_maskaddr_16 == 17)? _saxi_flag_17 : 
                            (axis_maskaddr_16 == 18)? _saxi_flag_18 : 
                            (axis_maskaddr_16 == 19)? _saxi_flag_19 : 
                            (axis_maskaddr_16 == 20)? _saxi_flag_20 : 
                            (axis_maskaddr_16 == 21)? _saxi_flag_21 : 
                            (axis_maskaddr_16 == 22)? _saxi_flag_22 : 
                            (axis_maskaddr_16 == 23)? _saxi_flag_23 : 
                            (axis_maskaddr_16 == 24)? _saxi_flag_24 : 
                            (axis_maskaddr_16 == 25)? _saxi_flag_25 : 
                            (axis_maskaddr_16 == 26)? _saxi_flag_26 : 
                            (axis_maskaddr_16 == 27)? _saxi_flag_27 : 
                            (axis_maskaddr_16 == 28)? _saxi_flag_28 : 
                            (axis_maskaddr_16 == 29)? _saxi_flag_29 : 
                            (axis_maskaddr_16 == 30)? _saxi_flag_30 : 
                            (axis_maskaddr_16 == 31)? _saxi_flag_31 : 
                            (axis_maskaddr_16 == 32)? _saxi_flag_32 : 
                            (axis_maskaddr_16 == 33)? _saxi_flag_33 : 
                            (axis_maskaddr_16 == 34)? _saxi_flag_34 : 
                            (axis_maskaddr_16 == 35)? _saxi_flag_35 : 
                            (axis_maskaddr_16 == 36)? _saxi_flag_36 : 'hx;
  wire signed [32-1:0] axislite_resetval_19;
  assign axislite_resetval_19 = (axis_maskaddr_16 == 0)? _saxi_resetval_0 : 
                                (axis_maskaddr_16 == 1)? _saxi_resetval_1 : 
                                (axis_maskaddr_16 == 2)? _saxi_resetval_2 : 
                                (axis_maskaddr_16 == 3)? _saxi_resetval_3 : 
                                (axis_maskaddr_16 == 4)? _saxi_resetval_4 : 
                                (axis_maskaddr_16 == 5)? _saxi_resetval_5 : 
                                (axis_maskaddr_16 == 6)? _saxi_resetval_6 : 
                                (axis_maskaddr_16 == 7)? _saxi_resetval_7 : 
                                (axis_maskaddr_16 == 8)? _saxi_resetval_8 : 
                                (axis_maskaddr_16 == 9)? _saxi_resetval_9 : 
                                (axis_maskaddr_16 == 10)? _saxi_resetval_10 : 
                                (axis_maskaddr_16 == 11)? _saxi_resetval_11 : 
                                (axis_maskaddr_16 == 12)? _saxi_resetval_12 : 
                                (axis_maskaddr_16 == 13)? _saxi_resetval_13 : 
                                (axis_maskaddr_16 == 14)? _saxi_resetval_14 : 
                                (axis_maskaddr_16 == 15)? _saxi_resetval_15 : 
                                (axis_maskaddr_16 == 16)? _saxi_resetval_16 : 
                                (axis_maskaddr_16 == 17)? _saxi_resetval_17 : 
                                (axis_maskaddr_16 == 18)? _saxi_resetval_18 : 
                                (axis_maskaddr_16 == 19)? _saxi_resetval_19 : 
                                (axis_maskaddr_16 == 20)? _saxi_resetval_20 : 
                                (axis_maskaddr_16 == 21)? _saxi_resetval_21 : 
                                (axis_maskaddr_16 == 22)? _saxi_resetval_22 : 
                                (axis_maskaddr_16 == 23)? _saxi_resetval_23 : 
                                (axis_maskaddr_16 == 24)? _saxi_resetval_24 : 
                                (axis_maskaddr_16 == 25)? _saxi_resetval_25 : 
                                (axis_maskaddr_16 == 26)? _saxi_resetval_26 : 
                                (axis_maskaddr_16 == 27)? _saxi_resetval_27 : 
                                (axis_maskaddr_16 == 28)? _saxi_resetval_28 : 
                                (axis_maskaddr_16 == 29)? _saxi_resetval_29 : 
                                (axis_maskaddr_16 == 30)? _saxi_resetval_30 : 
                                (axis_maskaddr_16 == 31)? _saxi_resetval_31 : 
                                (axis_maskaddr_16 == 32)? _saxi_resetval_32 : 
                                (axis_maskaddr_16 == 33)? _saxi_resetval_33 : 
                                (axis_maskaddr_16 == 34)? _saxi_resetval_34 : 
                                (axis_maskaddr_16 == 35)? _saxi_resetval_35 : 
                                (axis_maskaddr_16 == 36)? _saxi_resetval_36 : 'hx;
  reg _saxi_cond_0_1;
  assign saxi_wready = _saxi_register_fsm == 2;
  wire maxi_idle;
  assign maxi_idle = _maxi_write_idle & _maxi_read_idle;
  wire sw_rst_logic;
  assign sw_rst_logic = maxi_idle & _saxi_register_6;
  wire rst_logic;
  assign rst_logic = RESETN_inv_buf | sw_rst_logic;
  reg RST;
  reg _rst_logic_1;
  reg _rst_logic_2;
  wire signed [32-1:0] irq_20;
  assign irq_20 = _saxi_register_9 & _saxi_register_10;
  wire irq_busy;
  assign irq_busy = _saxi_register_5[0];
  reg irq_busy_edge_21;
  wire irq_busy_edge_22;
  assign irq_busy_edge_22 = irq_busy_edge_21 & !irq_busy;
  wire irq_extern;
  assign irq_extern = |_saxi_register_7;
  reg irq_extern_edge_23;
  wire irq_extern_edge_24;
  assign irq_extern_edge_24 = !irq_extern_edge_23 & irq_extern;
  wire [7-1:0] ram_w32_l128_id0_0_addr;
  wire [32-1:0] ram_w32_l128_id0_0_rdata;
  wire [32-1:0] ram_w32_l128_id0_0_wdata;
  wire ram_w32_l128_id0_0_wenable;
  wire ram_w32_l128_id0_0_enable;
  wire [7-1:0] ram_w32_l128_id0_1_addr;
  wire [32-1:0] ram_w32_l128_id0_1_rdata;
  wire [32-1:0] ram_w32_l128_id0_1_wdata;
  wire ram_w32_l128_id0_1_wenable;
  wire ram_w32_l128_id0_1_enable;

  ram_w32_l128_id0
  inst_ram_w32_l128_id0
  (
    .CLK(CLK),
    .ram_w32_l128_id0_0_addr(ram_w32_l128_id0_0_addr),
    .ram_w32_l128_id0_0_rdata(ram_w32_l128_id0_0_rdata),
    .ram_w32_l128_id0_0_wdata(ram_w32_l128_id0_0_wdata),
    .ram_w32_l128_id0_0_wenable(ram_w32_l128_id0_0_wenable),
    .ram_w32_l128_id0_0_enable(ram_w32_l128_id0_0_enable),
    .ram_w32_l128_id0_1_addr(ram_w32_l128_id0_1_addr),
    .ram_w32_l128_id0_1_rdata(ram_w32_l128_id0_1_rdata),
    .ram_w32_l128_id0_1_wdata(ram_w32_l128_id0_1_wdata),
    .ram_w32_l128_id0_1_wenable(ram_w32_l128_id0_1_wenable),
    .ram_w32_l128_id0_1_enable(ram_w32_l128_id0_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id1_0_addr;
  wire [32-1:0] ram_w32_l128_id1_0_rdata;
  wire [32-1:0] ram_w32_l128_id1_0_wdata;
  wire ram_w32_l128_id1_0_wenable;
  wire ram_w32_l128_id1_0_enable;
  wire [7-1:0] ram_w32_l128_id1_1_addr;
  wire [32-1:0] ram_w32_l128_id1_1_rdata;
  wire [32-1:0] ram_w32_l128_id1_1_wdata;
  wire ram_w32_l128_id1_1_wenable;
  wire ram_w32_l128_id1_1_enable;

  ram_w32_l128_id1
  inst_ram_w32_l128_id1
  (
    .CLK(CLK),
    .ram_w32_l128_id1_0_addr(ram_w32_l128_id1_0_addr),
    .ram_w32_l128_id1_0_rdata(ram_w32_l128_id1_0_rdata),
    .ram_w32_l128_id1_0_wdata(ram_w32_l128_id1_0_wdata),
    .ram_w32_l128_id1_0_wenable(ram_w32_l128_id1_0_wenable),
    .ram_w32_l128_id1_0_enable(ram_w32_l128_id1_0_enable),
    .ram_w32_l128_id1_1_addr(ram_w32_l128_id1_1_addr),
    .ram_w32_l128_id1_1_rdata(ram_w32_l128_id1_1_rdata),
    .ram_w32_l128_id1_1_wdata(ram_w32_l128_id1_1_wdata),
    .ram_w32_l128_id1_1_wenable(ram_w32_l128_id1_1_wenable),
    .ram_w32_l128_id1_1_enable(ram_w32_l128_id1_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id2_0_addr;
  wire [32-1:0] ram_w32_l128_id2_0_rdata;
  wire [32-1:0] ram_w32_l128_id2_0_wdata;
  wire ram_w32_l128_id2_0_wenable;
  wire ram_w32_l128_id2_0_enable;
  wire [7-1:0] ram_w32_l128_id2_1_addr;
  wire [32-1:0] ram_w32_l128_id2_1_rdata;
  wire [32-1:0] ram_w32_l128_id2_1_wdata;
  wire ram_w32_l128_id2_1_wenable;
  wire ram_w32_l128_id2_1_enable;
  assign ram_w32_l128_id2_0_wdata = 'hx;
  assign ram_w32_l128_id2_0_wenable = 0;

  ram_w32_l128_id2
  inst_ram_w32_l128_id2
  (
    .CLK(CLK),
    .ram_w32_l128_id2_0_addr(ram_w32_l128_id2_0_addr),
    .ram_w32_l128_id2_0_rdata(ram_w32_l128_id2_0_rdata),
    .ram_w32_l128_id2_0_wdata(ram_w32_l128_id2_0_wdata),
    .ram_w32_l128_id2_0_wenable(ram_w32_l128_id2_0_wenable),
    .ram_w32_l128_id2_0_enable(ram_w32_l128_id2_0_enable),
    .ram_w32_l128_id2_1_addr(ram_w32_l128_id2_1_addr),
    .ram_w32_l128_id2_1_rdata(ram_w32_l128_id2_1_rdata),
    .ram_w32_l128_id2_1_wdata(ram_w32_l128_id2_1_wdata),
    .ram_w32_l128_id2_1_wenable(ram_w32_l128_id2_1_wenable),
    .ram_w32_l128_id2_1_enable(ram_w32_l128_id2_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id3_0_addr;
  wire [32-1:0] ram_w32_l128_id3_0_rdata;
  wire [32-1:0] ram_w32_l128_id3_0_wdata;
  wire ram_w32_l128_id3_0_wenable;
  wire ram_w32_l128_id3_0_enable;
  wire [7-1:0] ram_w32_l128_id3_1_addr;
  wire [32-1:0] ram_w32_l128_id3_1_rdata;
  wire [32-1:0] ram_w32_l128_id3_1_wdata;
  wire ram_w32_l128_id3_1_wenable;
  wire ram_w32_l128_id3_1_enable;
  assign ram_w32_l128_id3_0_wdata = 'hx;
  assign ram_w32_l128_id3_0_wenable = 0;

  ram_w32_l128_id3
  inst_ram_w32_l128_id3
  (
    .CLK(CLK),
    .ram_w32_l128_id3_0_addr(ram_w32_l128_id3_0_addr),
    .ram_w32_l128_id3_0_rdata(ram_w32_l128_id3_0_rdata),
    .ram_w32_l128_id3_0_wdata(ram_w32_l128_id3_0_wdata),
    .ram_w32_l128_id3_0_wenable(ram_w32_l128_id3_0_wenable),
    .ram_w32_l128_id3_0_enable(ram_w32_l128_id3_0_enable),
    .ram_w32_l128_id3_1_addr(ram_w32_l128_id3_1_addr),
    .ram_w32_l128_id3_1_rdata(ram_w32_l128_id3_1_rdata),
    .ram_w32_l128_id3_1_wdata(ram_w32_l128_id3_1_wdata),
    .ram_w32_l128_id3_1_wenable(ram_w32_l128_id3_1_wenable),
    .ram_w32_l128_id3_1_enable(ram_w32_l128_id3_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id4_0_addr;
  wire [32-1:0] ram_w32_l128_id4_0_rdata;
  wire [32-1:0] ram_w32_l128_id4_0_wdata;
  wire ram_w32_l128_id4_0_wenable;
  wire ram_w32_l128_id4_0_enable;
  wire [7-1:0] ram_w32_l128_id4_1_addr;
  wire [32-1:0] ram_w32_l128_id4_1_rdata;
  wire [32-1:0] ram_w32_l128_id4_1_wdata;
  wire ram_w32_l128_id4_1_wenable;
  wire ram_w32_l128_id4_1_enable;
  assign ram_w32_l128_id4_0_wdata = 'hx;
  assign ram_w32_l128_id4_0_wenable = 0;

  ram_w32_l128_id4
  inst_ram_w32_l128_id4
  (
    .CLK(CLK),
    .ram_w32_l128_id4_0_addr(ram_w32_l128_id4_0_addr),
    .ram_w32_l128_id4_0_rdata(ram_w32_l128_id4_0_rdata),
    .ram_w32_l128_id4_0_wdata(ram_w32_l128_id4_0_wdata),
    .ram_w32_l128_id4_0_wenable(ram_w32_l128_id4_0_wenable),
    .ram_w32_l128_id4_0_enable(ram_w32_l128_id4_0_enable),
    .ram_w32_l128_id4_1_addr(ram_w32_l128_id4_1_addr),
    .ram_w32_l128_id4_1_rdata(ram_w32_l128_id4_1_rdata),
    .ram_w32_l128_id4_1_wdata(ram_w32_l128_id4_1_wdata),
    .ram_w32_l128_id4_1_wenable(ram_w32_l128_id4_1_wenable),
    .ram_w32_l128_id4_1_enable(ram_w32_l128_id4_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id5_0_addr;
  wire [32-1:0] ram_w32_l128_id5_0_rdata;
  wire [32-1:0] ram_w32_l128_id5_0_wdata;
  wire ram_w32_l128_id5_0_wenable;
  wire ram_w32_l128_id5_0_enable;
  wire [7-1:0] ram_w32_l128_id5_1_addr;
  wire [32-1:0] ram_w32_l128_id5_1_rdata;
  wire [32-1:0] ram_w32_l128_id5_1_wdata;
  wire ram_w32_l128_id5_1_wenable;
  wire ram_w32_l128_id5_1_enable;
  assign ram_w32_l128_id5_0_wdata = 'hx;
  assign ram_w32_l128_id5_0_wenable = 0;

  ram_w32_l128_id5
  inst_ram_w32_l128_id5
  (
    .CLK(CLK),
    .ram_w32_l128_id5_0_addr(ram_w32_l128_id5_0_addr),
    .ram_w32_l128_id5_0_rdata(ram_w32_l128_id5_0_rdata),
    .ram_w32_l128_id5_0_wdata(ram_w32_l128_id5_0_wdata),
    .ram_w32_l128_id5_0_wenable(ram_w32_l128_id5_0_wenable),
    .ram_w32_l128_id5_0_enable(ram_w32_l128_id5_0_enable),
    .ram_w32_l128_id5_1_addr(ram_w32_l128_id5_1_addr),
    .ram_w32_l128_id5_1_rdata(ram_w32_l128_id5_1_rdata),
    .ram_w32_l128_id5_1_wdata(ram_w32_l128_id5_1_wdata),
    .ram_w32_l128_id5_1_wenable(ram_w32_l128_id5_1_wenable),
    .ram_w32_l128_id5_1_enable(ram_w32_l128_id5_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id6_0_addr;
  wire [32-1:0] ram_w32_l128_id6_0_rdata;
  wire [32-1:0] ram_w32_l128_id6_0_wdata;
  wire ram_w32_l128_id6_0_wenable;
  wire ram_w32_l128_id6_0_enable;
  wire [7-1:0] ram_w32_l128_id6_1_addr;
  wire [32-1:0] ram_w32_l128_id6_1_rdata;
  wire [32-1:0] ram_w32_l128_id6_1_wdata;
  wire ram_w32_l128_id6_1_wenable;
  wire ram_w32_l128_id6_1_enable;
  assign ram_w32_l128_id6_0_wdata = 'hx;
  assign ram_w32_l128_id6_0_wenable = 0;

  ram_w32_l128_id6
  inst_ram_w32_l128_id6
  (
    .CLK(CLK),
    .ram_w32_l128_id6_0_addr(ram_w32_l128_id6_0_addr),
    .ram_w32_l128_id6_0_rdata(ram_w32_l128_id6_0_rdata),
    .ram_w32_l128_id6_0_wdata(ram_w32_l128_id6_0_wdata),
    .ram_w32_l128_id6_0_wenable(ram_w32_l128_id6_0_wenable),
    .ram_w32_l128_id6_0_enable(ram_w32_l128_id6_0_enable),
    .ram_w32_l128_id6_1_addr(ram_w32_l128_id6_1_addr),
    .ram_w32_l128_id6_1_rdata(ram_w32_l128_id6_1_rdata),
    .ram_w32_l128_id6_1_wdata(ram_w32_l128_id6_1_wdata),
    .ram_w32_l128_id6_1_wenable(ram_w32_l128_id6_1_wenable),
    .ram_w32_l128_id6_1_enable(ram_w32_l128_id6_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id7_0_addr;
  wire [32-1:0] ram_w32_l128_id7_0_rdata;
  wire [32-1:0] ram_w32_l128_id7_0_wdata;
  wire ram_w32_l128_id7_0_wenable;
  wire ram_w32_l128_id7_0_enable;
  wire [7-1:0] ram_w32_l128_id7_1_addr;
  wire [32-1:0] ram_w32_l128_id7_1_rdata;
  wire [32-1:0] ram_w32_l128_id7_1_wdata;
  wire ram_w32_l128_id7_1_wenable;
  wire ram_w32_l128_id7_1_enable;
  assign ram_w32_l128_id7_0_wdata = 'hx;
  assign ram_w32_l128_id7_0_wenable = 0;

  ram_w32_l128_id7
  inst_ram_w32_l128_id7
  (
    .CLK(CLK),
    .ram_w32_l128_id7_0_addr(ram_w32_l128_id7_0_addr),
    .ram_w32_l128_id7_0_rdata(ram_w32_l128_id7_0_rdata),
    .ram_w32_l128_id7_0_wdata(ram_w32_l128_id7_0_wdata),
    .ram_w32_l128_id7_0_wenable(ram_w32_l128_id7_0_wenable),
    .ram_w32_l128_id7_0_enable(ram_w32_l128_id7_0_enable),
    .ram_w32_l128_id7_1_addr(ram_w32_l128_id7_1_addr),
    .ram_w32_l128_id7_1_rdata(ram_w32_l128_id7_1_rdata),
    .ram_w32_l128_id7_1_wdata(ram_w32_l128_id7_1_wdata),
    .ram_w32_l128_id7_1_wenable(ram_w32_l128_id7_1_wenable),
    .ram_w32_l128_id7_1_enable(ram_w32_l128_id7_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id8_0_addr;
  wire [32-1:0] ram_w32_l128_id8_0_rdata;
  wire [32-1:0] ram_w32_l128_id8_0_wdata;
  wire ram_w32_l128_id8_0_wenable;
  wire ram_w32_l128_id8_0_enable;
  wire [7-1:0] ram_w32_l128_id8_1_addr;
  wire [32-1:0] ram_w32_l128_id8_1_rdata;
  wire [32-1:0] ram_w32_l128_id8_1_wdata;
  wire ram_w32_l128_id8_1_wenable;
  wire ram_w32_l128_id8_1_enable;
  assign ram_w32_l128_id8_0_wdata = 'hx;
  assign ram_w32_l128_id8_0_wenable = 0;

  ram_w32_l128_id8
  inst_ram_w32_l128_id8
  (
    .CLK(CLK),
    .ram_w32_l128_id8_0_addr(ram_w32_l128_id8_0_addr),
    .ram_w32_l128_id8_0_rdata(ram_w32_l128_id8_0_rdata),
    .ram_w32_l128_id8_0_wdata(ram_w32_l128_id8_0_wdata),
    .ram_w32_l128_id8_0_wenable(ram_w32_l128_id8_0_wenable),
    .ram_w32_l128_id8_0_enable(ram_w32_l128_id8_0_enable),
    .ram_w32_l128_id8_1_addr(ram_w32_l128_id8_1_addr),
    .ram_w32_l128_id8_1_rdata(ram_w32_l128_id8_1_rdata),
    .ram_w32_l128_id8_1_wdata(ram_w32_l128_id8_1_wdata),
    .ram_w32_l128_id8_1_wenable(ram_w32_l128_id8_1_wenable),
    .ram_w32_l128_id8_1_enable(ram_w32_l128_id8_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id9_0_addr;
  wire [32-1:0] ram_w32_l128_id9_0_rdata;
  wire [32-1:0] ram_w32_l128_id9_0_wdata;
  wire ram_w32_l128_id9_0_wenable;
  wire ram_w32_l128_id9_0_enable;
  wire [7-1:0] ram_w32_l128_id9_1_addr;
  wire [32-1:0] ram_w32_l128_id9_1_rdata;
  wire [32-1:0] ram_w32_l128_id9_1_wdata;
  wire ram_w32_l128_id9_1_wenable;
  wire ram_w32_l128_id9_1_enable;
  assign ram_w32_l128_id9_0_wdata = 'hx;
  assign ram_w32_l128_id9_0_wenable = 0;

  ram_w32_l128_id9
  inst_ram_w32_l128_id9
  (
    .CLK(CLK),
    .ram_w32_l128_id9_0_addr(ram_w32_l128_id9_0_addr),
    .ram_w32_l128_id9_0_rdata(ram_w32_l128_id9_0_rdata),
    .ram_w32_l128_id9_0_wdata(ram_w32_l128_id9_0_wdata),
    .ram_w32_l128_id9_0_wenable(ram_w32_l128_id9_0_wenable),
    .ram_w32_l128_id9_0_enable(ram_w32_l128_id9_0_enable),
    .ram_w32_l128_id9_1_addr(ram_w32_l128_id9_1_addr),
    .ram_w32_l128_id9_1_rdata(ram_w32_l128_id9_1_rdata),
    .ram_w32_l128_id9_1_wdata(ram_w32_l128_id9_1_wdata),
    .ram_w32_l128_id9_1_wenable(ram_w32_l128_id9_1_wenable),
    .ram_w32_l128_id9_1_enable(ram_w32_l128_id9_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id10_0_addr;
  wire [32-1:0] ram_w32_l128_id10_0_rdata;
  wire [32-1:0] ram_w32_l128_id10_0_wdata;
  wire ram_w32_l128_id10_0_wenable;
  wire ram_w32_l128_id10_0_enable;
  wire [7-1:0] ram_w32_l128_id10_1_addr;
  wire [32-1:0] ram_w32_l128_id10_1_rdata;
  wire [32-1:0] ram_w32_l128_id10_1_wdata;
  wire ram_w32_l128_id10_1_wenable;
  wire ram_w32_l128_id10_1_enable;
  assign ram_w32_l128_id10_0_wdata = 'hx;
  assign ram_w32_l128_id10_0_wenable = 0;

  ram_w32_l128_id10
  inst_ram_w32_l128_id10
  (
    .CLK(CLK),
    .ram_w32_l128_id10_0_addr(ram_w32_l128_id10_0_addr),
    .ram_w32_l128_id10_0_rdata(ram_w32_l128_id10_0_rdata),
    .ram_w32_l128_id10_0_wdata(ram_w32_l128_id10_0_wdata),
    .ram_w32_l128_id10_0_wenable(ram_w32_l128_id10_0_wenable),
    .ram_w32_l128_id10_0_enable(ram_w32_l128_id10_0_enable),
    .ram_w32_l128_id10_1_addr(ram_w32_l128_id10_1_addr),
    .ram_w32_l128_id10_1_rdata(ram_w32_l128_id10_1_rdata),
    .ram_w32_l128_id10_1_wdata(ram_w32_l128_id10_1_wdata),
    .ram_w32_l128_id10_1_wenable(ram_w32_l128_id10_1_wenable),
    .ram_w32_l128_id10_1_enable(ram_w32_l128_id10_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id11_0_addr;
  wire [32-1:0] ram_w32_l128_id11_0_rdata;
  wire [32-1:0] ram_w32_l128_id11_0_wdata;
  wire ram_w32_l128_id11_0_wenable;
  wire ram_w32_l128_id11_0_enable;
  wire [7-1:0] ram_w32_l128_id11_1_addr;
  wire [32-1:0] ram_w32_l128_id11_1_rdata;
  wire [32-1:0] ram_w32_l128_id11_1_wdata;
  wire ram_w32_l128_id11_1_wenable;
  wire ram_w32_l128_id11_1_enable;
  assign ram_w32_l128_id11_0_wdata = 'hx;
  assign ram_w32_l128_id11_0_wenable = 0;

  ram_w32_l128_id11
  inst_ram_w32_l128_id11
  (
    .CLK(CLK),
    .ram_w32_l128_id11_0_addr(ram_w32_l128_id11_0_addr),
    .ram_w32_l128_id11_0_rdata(ram_w32_l128_id11_0_rdata),
    .ram_w32_l128_id11_0_wdata(ram_w32_l128_id11_0_wdata),
    .ram_w32_l128_id11_0_wenable(ram_w32_l128_id11_0_wenable),
    .ram_w32_l128_id11_0_enable(ram_w32_l128_id11_0_enable),
    .ram_w32_l128_id11_1_addr(ram_w32_l128_id11_1_addr),
    .ram_w32_l128_id11_1_rdata(ram_w32_l128_id11_1_rdata),
    .ram_w32_l128_id11_1_wdata(ram_w32_l128_id11_1_wdata),
    .ram_w32_l128_id11_1_wenable(ram_w32_l128_id11_1_wenable),
    .ram_w32_l128_id11_1_enable(ram_w32_l128_id11_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id12_0_addr;
  wire [32-1:0] ram_w32_l128_id12_0_rdata;
  wire [32-1:0] ram_w32_l128_id12_0_wdata;
  wire ram_w32_l128_id12_0_wenable;
  wire ram_w32_l128_id12_0_enable;
  wire [7-1:0] ram_w32_l128_id12_1_addr;
  wire [32-1:0] ram_w32_l128_id12_1_rdata;
  wire [32-1:0] ram_w32_l128_id12_1_wdata;
  wire ram_w32_l128_id12_1_wenable;
  wire ram_w32_l128_id12_1_enable;
  assign ram_w32_l128_id12_0_wdata = 'hx;
  assign ram_w32_l128_id12_0_wenable = 0;

  ram_w32_l128_id12
  inst_ram_w32_l128_id12
  (
    .CLK(CLK),
    .ram_w32_l128_id12_0_addr(ram_w32_l128_id12_0_addr),
    .ram_w32_l128_id12_0_rdata(ram_w32_l128_id12_0_rdata),
    .ram_w32_l128_id12_0_wdata(ram_w32_l128_id12_0_wdata),
    .ram_w32_l128_id12_0_wenable(ram_w32_l128_id12_0_wenable),
    .ram_w32_l128_id12_0_enable(ram_w32_l128_id12_0_enable),
    .ram_w32_l128_id12_1_addr(ram_w32_l128_id12_1_addr),
    .ram_w32_l128_id12_1_rdata(ram_w32_l128_id12_1_rdata),
    .ram_w32_l128_id12_1_wdata(ram_w32_l128_id12_1_wdata),
    .ram_w32_l128_id12_1_wenable(ram_w32_l128_id12_1_wenable),
    .ram_w32_l128_id12_1_enable(ram_w32_l128_id12_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id13_0_addr;
  wire [32-1:0] ram_w32_l128_id13_0_rdata;
  wire [32-1:0] ram_w32_l128_id13_0_wdata;
  wire ram_w32_l128_id13_0_wenable;
  wire ram_w32_l128_id13_0_enable;
  wire [7-1:0] ram_w32_l128_id13_1_addr;
  wire [32-1:0] ram_w32_l128_id13_1_rdata;
  wire [32-1:0] ram_w32_l128_id13_1_wdata;
  wire ram_w32_l128_id13_1_wenable;
  wire ram_w32_l128_id13_1_enable;
  assign ram_w32_l128_id13_0_wdata = 'hx;
  assign ram_w32_l128_id13_0_wenable = 0;

  ram_w32_l128_id13
  inst_ram_w32_l128_id13
  (
    .CLK(CLK),
    .ram_w32_l128_id13_0_addr(ram_w32_l128_id13_0_addr),
    .ram_w32_l128_id13_0_rdata(ram_w32_l128_id13_0_rdata),
    .ram_w32_l128_id13_0_wdata(ram_w32_l128_id13_0_wdata),
    .ram_w32_l128_id13_0_wenable(ram_w32_l128_id13_0_wenable),
    .ram_w32_l128_id13_0_enable(ram_w32_l128_id13_0_enable),
    .ram_w32_l128_id13_1_addr(ram_w32_l128_id13_1_addr),
    .ram_w32_l128_id13_1_rdata(ram_w32_l128_id13_1_rdata),
    .ram_w32_l128_id13_1_wdata(ram_w32_l128_id13_1_wdata),
    .ram_w32_l128_id13_1_wenable(ram_w32_l128_id13_1_wenable),
    .ram_w32_l128_id13_1_enable(ram_w32_l128_id13_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id14_0_addr;
  wire [32-1:0] ram_w32_l128_id14_0_rdata;
  wire [32-1:0] ram_w32_l128_id14_0_wdata;
  wire ram_w32_l128_id14_0_wenable;
  wire ram_w32_l128_id14_0_enable;
  wire [7-1:0] ram_w32_l128_id14_1_addr;
  wire [32-1:0] ram_w32_l128_id14_1_rdata;
  wire [32-1:0] ram_w32_l128_id14_1_wdata;
  wire ram_w32_l128_id14_1_wenable;
  wire ram_w32_l128_id14_1_enable;
  assign ram_w32_l128_id14_0_wdata = 'hx;
  assign ram_w32_l128_id14_0_wenable = 0;

  ram_w32_l128_id14
  inst_ram_w32_l128_id14
  (
    .CLK(CLK),
    .ram_w32_l128_id14_0_addr(ram_w32_l128_id14_0_addr),
    .ram_w32_l128_id14_0_rdata(ram_w32_l128_id14_0_rdata),
    .ram_w32_l128_id14_0_wdata(ram_w32_l128_id14_0_wdata),
    .ram_w32_l128_id14_0_wenable(ram_w32_l128_id14_0_wenable),
    .ram_w32_l128_id14_0_enable(ram_w32_l128_id14_0_enable),
    .ram_w32_l128_id14_1_addr(ram_w32_l128_id14_1_addr),
    .ram_w32_l128_id14_1_rdata(ram_w32_l128_id14_1_rdata),
    .ram_w32_l128_id14_1_wdata(ram_w32_l128_id14_1_wdata),
    .ram_w32_l128_id14_1_wenable(ram_w32_l128_id14_1_wenable),
    .ram_w32_l128_id14_1_enable(ram_w32_l128_id14_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id15_0_addr;
  wire [32-1:0] ram_w32_l128_id15_0_rdata;
  wire [32-1:0] ram_w32_l128_id15_0_wdata;
  wire ram_w32_l128_id15_0_wenable;
  wire ram_w32_l128_id15_0_enable;
  wire [7-1:0] ram_w32_l128_id15_1_addr;
  wire [32-1:0] ram_w32_l128_id15_1_rdata;
  wire [32-1:0] ram_w32_l128_id15_1_wdata;
  wire ram_w32_l128_id15_1_wenable;
  wire ram_w32_l128_id15_1_enable;
  assign ram_w32_l128_id15_0_wdata = 'hx;
  assign ram_w32_l128_id15_0_wenable = 0;

  ram_w32_l128_id15
  inst_ram_w32_l128_id15
  (
    .CLK(CLK),
    .ram_w32_l128_id15_0_addr(ram_w32_l128_id15_0_addr),
    .ram_w32_l128_id15_0_rdata(ram_w32_l128_id15_0_rdata),
    .ram_w32_l128_id15_0_wdata(ram_w32_l128_id15_0_wdata),
    .ram_w32_l128_id15_0_wenable(ram_w32_l128_id15_0_wenable),
    .ram_w32_l128_id15_0_enable(ram_w32_l128_id15_0_enable),
    .ram_w32_l128_id15_1_addr(ram_w32_l128_id15_1_addr),
    .ram_w32_l128_id15_1_rdata(ram_w32_l128_id15_1_rdata),
    .ram_w32_l128_id15_1_wdata(ram_w32_l128_id15_1_wdata),
    .ram_w32_l128_id15_1_wenable(ram_w32_l128_id15_1_wenable),
    .ram_w32_l128_id15_1_enable(ram_w32_l128_id15_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id16_0_addr;
  wire [32-1:0] ram_w32_l128_id16_0_rdata;
  wire [32-1:0] ram_w32_l128_id16_0_wdata;
  wire ram_w32_l128_id16_0_wenable;
  wire ram_w32_l128_id16_0_enable;
  wire [7-1:0] ram_w32_l128_id16_1_addr;
  wire [32-1:0] ram_w32_l128_id16_1_rdata;
  wire [32-1:0] ram_w32_l128_id16_1_wdata;
  wire ram_w32_l128_id16_1_wenable;
  wire ram_w32_l128_id16_1_enable;
  assign ram_w32_l128_id16_0_wdata = 'hx;
  assign ram_w32_l128_id16_0_wenable = 0;

  ram_w32_l128_id16
  inst_ram_w32_l128_id16
  (
    .CLK(CLK),
    .ram_w32_l128_id16_0_addr(ram_w32_l128_id16_0_addr),
    .ram_w32_l128_id16_0_rdata(ram_w32_l128_id16_0_rdata),
    .ram_w32_l128_id16_0_wdata(ram_w32_l128_id16_0_wdata),
    .ram_w32_l128_id16_0_wenable(ram_w32_l128_id16_0_wenable),
    .ram_w32_l128_id16_0_enable(ram_w32_l128_id16_0_enable),
    .ram_w32_l128_id16_1_addr(ram_w32_l128_id16_1_addr),
    .ram_w32_l128_id16_1_rdata(ram_w32_l128_id16_1_rdata),
    .ram_w32_l128_id16_1_wdata(ram_w32_l128_id16_1_wdata),
    .ram_w32_l128_id16_1_wenable(ram_w32_l128_id16_1_wenable),
    .ram_w32_l128_id16_1_enable(ram_w32_l128_id16_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id17_0_addr;
  wire [32-1:0] ram_w32_l128_id17_0_rdata;
  wire [32-1:0] ram_w32_l128_id17_0_wdata;
  wire ram_w32_l128_id17_0_wenable;
  wire ram_w32_l128_id17_0_enable;
  wire [7-1:0] ram_w32_l128_id17_1_addr;
  wire [32-1:0] ram_w32_l128_id17_1_rdata;
  wire [32-1:0] ram_w32_l128_id17_1_wdata;
  wire ram_w32_l128_id17_1_wenable;
  wire ram_w32_l128_id17_1_enable;
  assign ram_w32_l128_id17_0_wdata = 'hx;
  assign ram_w32_l128_id17_0_wenable = 0;

  ram_w32_l128_id17
  inst_ram_w32_l128_id17
  (
    .CLK(CLK),
    .ram_w32_l128_id17_0_addr(ram_w32_l128_id17_0_addr),
    .ram_w32_l128_id17_0_rdata(ram_w32_l128_id17_0_rdata),
    .ram_w32_l128_id17_0_wdata(ram_w32_l128_id17_0_wdata),
    .ram_w32_l128_id17_0_wenable(ram_w32_l128_id17_0_wenable),
    .ram_w32_l128_id17_0_enable(ram_w32_l128_id17_0_enable),
    .ram_w32_l128_id17_1_addr(ram_w32_l128_id17_1_addr),
    .ram_w32_l128_id17_1_rdata(ram_w32_l128_id17_1_rdata),
    .ram_w32_l128_id17_1_wdata(ram_w32_l128_id17_1_wdata),
    .ram_w32_l128_id17_1_wenable(ram_w32_l128_id17_1_wenable),
    .ram_w32_l128_id17_1_enable(ram_w32_l128_id17_1_enable)
  );

  wire [7-1:0] ram_w32_l128_id18_0_addr;
  wire [32-1:0] ram_w32_l128_id18_0_rdata;
  wire [32-1:0] ram_w32_l128_id18_0_wdata;
  wire ram_w32_l128_id18_0_wenable;
  wire ram_w32_l128_id18_0_enable;
  wire [7-1:0] ram_w32_l128_id18_1_addr;
  wire [32-1:0] ram_w32_l128_id18_1_rdata;
  wire [32-1:0] ram_w32_l128_id18_1_wdata;
  wire ram_w32_l128_id18_1_wenable;
  wire ram_w32_l128_id18_1_enable;
  assign ram_w32_l128_id18_0_wdata = 'hx;
  assign ram_w32_l128_id18_0_wenable = 0;

  ram_w32_l128_id18
  inst_ram_w32_l128_id18
  (
    .CLK(CLK),
    .ram_w32_l128_id18_0_addr(ram_w32_l128_id18_0_addr),
    .ram_w32_l128_id18_0_rdata(ram_w32_l128_id18_0_rdata),
    .ram_w32_l128_id18_0_wdata(ram_w32_l128_id18_0_wdata),
    .ram_w32_l128_id18_0_wenable(ram_w32_l128_id18_0_wenable),
    .ram_w32_l128_id18_0_enable(ram_w32_l128_id18_0_enable),
    .ram_w32_l128_id18_1_addr(ram_w32_l128_id18_1_addr),
    .ram_w32_l128_id18_1_rdata(ram_w32_l128_id18_1_rdata),
    .ram_w32_l128_id18_1_wdata(ram_w32_l128_id18_1_wdata),
    .ram_w32_l128_id18_1_wenable(ram_w32_l128_id18_1_wenable),
    .ram_w32_l128_id18_1_enable(ram_w32_l128_id18_1_enable)
  );

  wire [3-1:0] cparam_conv2d_2_act_num_col;
  wire [3-1:0] cparam_conv2d_2_act_num_row;
  wire [3-1:0] cparam_conv2d_2_filter_num_och;
  wire [1-1:0] cparam_conv2d_2_bias_scala;
  wire [1-1:0] cparam_conv2d_2_bias_num;
  wire [1-1:0] cparam_conv2d_2_scale_scala;
  wire [1-1:0] cparam_conv2d_2_scale_num;
  wire [1-1:0] cparam_conv2d_2_vshamt_mul_scala;
  wire [1-1:0] cparam_conv2d_2_vshamt_mul_num;
  wire [1-1:0] cparam_conv2d_2_vshamt_sum_scala;
  wire [1-1:0] cparam_conv2d_2_vshamt_sum_num;
  wire [1-1:0] cparam_conv2d_2_vshamt_out_scala;
  wire [1-1:0] cparam_conv2d_2_vshamt_out_num;
  wire [1-1:0] cparam_conv2d_2_cshamt_mul_value;
  wire [1-1:0] cparam_conv2d_2_cshamt_sum_value;
  wire [1-1:0] cparam_conv2d_2_cshamt_out_value;
  wire [1-1:0] cparam_conv2d_2_act_func_index;
  wire [3-1:0] cparam_conv2d_2_out_num_col;
  wire [3-1:0] cparam_conv2d_2_out_num_row;
  wire [1-1:0] cparam_conv2d_2_pad_col_left;
  wire [1-1:0] cparam_conv2d_2_pad_row_top;
  wire [3-1:0] cparam_conv2d_2_max_col_count;
  wire [3-1:0] cparam_conv2d_2_max_row_count;
  wire [1-1:0] cparam_conv2d_2_max_bat_count;
  wire [2-1:0] cparam_conv2d_2_max_och_count;
  wire [3-1:0] cparam_conv2d_2_och_count_step;
  wire [1-1:0] cparam_conv2d_2_dma_flag_conds_0;
  wire [1-1:0] cparam_conv2d_2_dma_flag_conds_1;
  wire [1-1:0] cparam_conv2d_2_dma_flag_conds_2;
  wire signed [32-1:0] cparam_conv2d_2_act_offset_values_0;
  wire signed [32-1:0] cparam_conv2d_2_act_offset_values_1;
  wire signed [32-1:0] cparam_conv2d_2_act_offset_values_2;
  wire [9-1:0] cparam_conv2d_2_act_row_step;
  wire [12-1:0] cparam_conv2d_2_act_bat_step;
  wire [7-1:0] cparam_conv2d_2_act_read_size;
  wire [4-1:0] cparam_conv2d_2_act_read_block;
  wire [6-1:0] cparam_conv2d_2_act_read_step;
  wire [12-1:0] cparam_conv2d_2_filter_base_step;
  wire [10-1:0] cparam_conv2d_2_filter_read_size;
  wire [4-1:0] cparam_conv2d_2_filter_read_block;
  wire [6-1:0] cparam_conv2d_2_filter_read_step;
  wire [1-1:0] cparam_conv2d_2_out_offset_values_0;
  wire [5-1:0] cparam_conv2d_2_out_col_step;
  wire [8-1:0] cparam_conv2d_2_out_row_step;
  wire [11-1:0] cparam_conv2d_2_out_bat_step;
  wire [5-1:0] cparam_conv2d_2_out_och_step;
  wire [3-1:0] cparam_conv2d_2_out_write_size;
  wire [2-1:0] cparam_conv2d_2_out_write_size_res;
  wire [1-1:0] cparam_conv2d_2_out_write_block;
  wire [1-1:0] cparam_conv2d_2_keep_filter;
  wire [1-1:0] cparam_conv2d_2_keep_input;
  wire [1-1:0] cparam_conv2d_2_data_stationary;
  wire [3-1:0] cparam_conv2d_2_stream_num_ops;
  wire [2-1:0] cparam_conv2d_2_stream_num_ops_res;
  wire [3-1:0] cparam_conv2d_2_stream_num_ops_par;
  wire [2-1:0] cparam_conv2d_2_stream_num_ops_res_par;
  wire [4-1:0] cparam_conv2d_2_stream_reduce_size;
  wire [4-1:0] cparam_conv2d_2_stream_aligned_reduce_size;
  wire [1-1:0] cparam_conv2d_2_stream_omit_mask;
  wire [2-1:0] cparam_conv2d_2_col_select_initval;
  wire [1-1:0] cparam_conv2d_2_stride_col_par_col;
  wire [1-1:0] cparam_conv2d_2_stride_row_par_row;
  wire [1-1:0] cparam_conv2d_2_stride_col_mod_filter_num;
  wire [2-1:0] cparam_conv2d_2_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_8;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_9;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_10;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_11;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_12;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_13;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_14;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_15;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_16;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_17;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_18;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_19;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_20;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_21;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_22;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_23;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_24;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_25;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_conds_26;
  wire [1-1:0] cparam_conv2d_2_inc_act_laddr_small;
  wire [4-1:0] cparam_conv2d_2_inc_act_laddr_large;
  wire [3-1:0] cparam_conv2d_2_inc_out_laddr_col;
  wire [1-1:0] cparam_conv2d_2_stream_act_local_small_offset;
  wire signed [5-1:0] cparam_conv2d_2_stream_act_local_large_offset;
  wire [1-1:0] cparam_conv2d_2_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_conv2d_2_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_conv2d_2_stream_act_local_small_flags_2;
  wire [1-1:0] cparam_conv2d_2_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_conv2d_2_stream_act_local_large_flags_1;
  wire [1-1:0] cparam_conv2d_2_stream_act_local_large_flags_2;
  wire [1-1:0] cparam_conv2d_2_inc_sync_out;
  wire [1-1:0] cparam_conv2d_2_inc_sync_out_res;
  assign cparam_conv2d_2_act_num_col = 7;
  assign cparam_conv2d_2_act_num_row = 7;
  assign cparam_conv2d_2_filter_num_och = 7;
  assign cparam_conv2d_2_bias_scala = 0;
  assign cparam_conv2d_2_bias_num = 0;
  assign cparam_conv2d_2_scale_scala = 0;
  assign cparam_conv2d_2_scale_num = 0;
  assign cparam_conv2d_2_vshamt_mul_scala = 0;
  assign cparam_conv2d_2_vshamt_mul_num = 0;
  assign cparam_conv2d_2_vshamt_sum_scala = 0;
  assign cparam_conv2d_2_vshamt_sum_num = 0;
  assign cparam_conv2d_2_vshamt_out_scala = 0;
  assign cparam_conv2d_2_vshamt_out_num = 0;
  assign cparam_conv2d_2_cshamt_mul_value = 0;
  assign cparam_conv2d_2_cshamt_sum_value = 0;
  assign cparam_conv2d_2_cshamt_out_value = 0;
  assign cparam_conv2d_2_act_func_index = 0;
  assign cparam_conv2d_2_out_num_col = 7;
  assign cparam_conv2d_2_out_num_row = 7;
  assign cparam_conv2d_2_pad_col_left = 1;
  assign cparam_conv2d_2_pad_row_top = 1;
  assign cparam_conv2d_2_max_col_count = 6;
  assign cparam_conv2d_2_max_row_count = 6;
  assign cparam_conv2d_2_max_bat_count = 0;
  assign cparam_conv2d_2_max_och_count = 3;
  assign cparam_conv2d_2_och_count_step = 4;
  assign cparam_conv2d_2_dma_flag_conds_0 = 1;
  assign cparam_conv2d_2_dma_flag_conds_1 = 0;
  assign cparam_conv2d_2_dma_flag_conds_2 = 0;
  assign cparam_conv2d_2_act_offset_values_0 = -420;
  assign cparam_conv2d_2_act_offset_values_1 = 0;
  assign cparam_conv2d_2_act_offset_values_2 = 420;
  assign cparam_conv2d_2_act_row_step = 420;
  assign cparam_conv2d_2_act_bat_step = 2940;
  assign cparam_conv2d_2_act_read_size = 105;
  assign cparam_conv2d_2_act_read_block = 15;
  assign cparam_conv2d_2_act_read_step = 45;
  assign cparam_conv2d_2_filter_base_step = 2160;
  assign cparam_conv2d_2_filter_read_size = 540;
  assign cparam_conv2d_2_filter_read_block = 15;
  assign cparam_conv2d_2_filter_read_step = 60;
  assign cparam_conv2d_2_out_offset_values_0 = 0;
  assign cparam_conv2d_2_out_col_step = 28;
  assign cparam_conv2d_2_out_row_step = 196;
  assign cparam_conv2d_2_out_bat_step = 1372;
  assign cparam_conv2d_2_out_och_step = 16;
  assign cparam_conv2d_2_out_write_size = 4;
  assign cparam_conv2d_2_out_write_size_res = 3;
  assign cparam_conv2d_2_out_write_block = 0;
  assign cparam_conv2d_2_keep_filter = 0;
  assign cparam_conv2d_2_keep_input = 0;
  assign cparam_conv2d_2_data_stationary = 0;
  assign cparam_conv2d_2_stream_num_ops = 4;
  assign cparam_conv2d_2_stream_num_ops_res = 3;
  assign cparam_conv2d_2_stream_num_ops_par = 4;
  assign cparam_conv2d_2_stream_num_ops_res_par = 3;
  assign cparam_conv2d_2_stream_reduce_size = 15;
  assign cparam_conv2d_2_stream_aligned_reduce_size = 15;
  assign cparam_conv2d_2_stream_omit_mask = 0;
  assign cparam_conv2d_2_col_select_initval = 2;
  assign cparam_conv2d_2_stride_col_par_col = 1;
  assign cparam_conv2d_2_stride_row_par_row = 1;
  assign cparam_conv2d_2_stride_col_mod_filter_num = 1;
  assign cparam_conv2d_2_filter_num_col_minus_stride_col_mod = 2;
  assign cparam_conv2d_2_inc_act_laddr_conds_0 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_1 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_2 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_3 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_4 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_5 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_6 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_7 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_8 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_9 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_10 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_11 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_12 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_13 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_14 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_15 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_16 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_17 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_18 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_19 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_20 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_21 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_22 = 1;
  assign cparam_conv2d_2_inc_act_laddr_conds_23 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_24 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_25 = 0;
  assign cparam_conv2d_2_inc_act_laddr_conds_26 = 1;
  assign cparam_conv2d_2_inc_act_laddr_small = 0;
  assign cparam_conv2d_2_inc_act_laddr_large = 15;
  assign cparam_conv2d_2_inc_out_laddr_col = 7;
  assign cparam_conv2d_2_stream_act_local_small_offset = 0;
  assign cparam_conv2d_2_stream_act_local_large_offset = -15;
  assign cparam_conv2d_2_stream_act_local_small_flags_0 = 0;
  assign cparam_conv2d_2_stream_act_local_small_flags_1 = 0;
  assign cparam_conv2d_2_stream_act_local_small_flags_2 = 1;
  assign cparam_conv2d_2_stream_act_local_large_flags_0 = 0;
  assign cparam_conv2d_2_stream_act_local_large_flags_1 = 0;
  assign cparam_conv2d_2_stream_act_local_large_flags_2 = 1;
  assign cparam_conv2d_2_inc_sync_out = 1;
  assign cparam_conv2d_2_inc_sync_out_res = 0;
  wire [3-1:0] cparam_celu_3_dma_size;
  wire [6-1:0] cparam_celu_3_num_comp;
  wire [5-1:0] cparam_celu_3_addr_inc;
  wire [11-1:0] cparam_celu_3_arg_addr_incs_0;
  wire [8-1:0] cparam_celu_3_arg_addr_incs_1;
  wire [5-1:0] cparam_celu_3_arg_addr_incs_2;
  wire [1-1:0] cparam_celu_3_arg_addr_incs_3;
  wire [1-1:0] cparam_celu_3_arg_trip_sizes_0;
  wire [3-1:0] cparam_celu_3_arg_trip_sizes_1;
  wire [3-1:0] cparam_celu_3_arg_trip_sizes_2;
  wire [3-1:0] cparam_celu_3_arg_trip_sizes_3;
  wire [1-1:0] cparam_celu_3_arg_repeat_sizes_0;
  wire [1-1:0] cparam_celu_3_arg_repeat_sizes_1;
  wire [1-1:0] cparam_celu_3_arg_repeat_sizes_2;
  wire [1-1:0] cparam_celu_3_arg_repeat_sizes_3;
  wire [1-1:0] cparam_celu_3_arg_omit_dmas_0;
  wire [1-1:0] cparam_celu_3_arg_stride_zeros_0;
  wire [6-1:0] cparam_celu_3_local_0_features_scale_cparam;
  wire [1-1:0] cparam_celu_3_local_0_features_shamt_cparam;
  assign cparam_celu_3_dma_size = 7;
  assign cparam_celu_3_num_comp = 49;
  assign cparam_celu_3_addr_inc = 28;
  assign cparam_celu_3_arg_addr_incs_0 = 1372;
  assign cparam_celu_3_arg_addr_incs_1 = 196;
  assign cparam_celu_3_arg_addr_incs_2 = 28;
  assign cparam_celu_3_arg_addr_incs_3 = 0;
  assign cparam_celu_3_arg_trip_sizes_0 = 1;
  assign cparam_celu_3_arg_trip_sizes_1 = 7;
  assign cparam_celu_3_arg_trip_sizes_2 = 7;
  assign cparam_celu_3_arg_trip_sizes_3 = 7;
  assign cparam_celu_3_arg_repeat_sizes_0 = 1;
  assign cparam_celu_3_arg_repeat_sizes_1 = 1;
  assign cparam_celu_3_arg_repeat_sizes_2 = 1;
  assign cparam_celu_3_arg_repeat_sizes_3 = 1;
  assign cparam_celu_3_arg_omit_dmas_0 = 0;
  assign cparam_celu_3_arg_stride_zeros_0 = 0;
  assign cparam_celu_3_local_0_features_scale_cparam = 43;
  assign cparam_celu_3_local_0_features_shamt_cparam = 0;
  reg _acc_0_stream_ivalid;
  wire _acc_0_stream_oready;
  wire _acc_0_stream_internal_oready;
  assign _acc_0_stream_internal_oready = 1;
  reg [32-1:0] _acc_0_fsm;
  localparam _acc_0_fsm_init = 0;
  wire _acc_0_run_flag;
  assign _acc_0_run_flag = 0;
  reg _acc_0_source_start;
  wire _acc_0_source_stop;
  reg _acc_0_source_busy;
  wire _acc_0_sink_start;
  wire _acc_0_sink_stop;
  wire _acc_0_sink_busy;
  wire _acc_0_busy;
  reg _acc_0_busy_reg;
  wire _acc_0_is_root;
  reg _acc_0_x_idle;
  reg [33-1:0] _acc_0_x_source_count;
  reg [5-1:0] _acc_0_x_source_mode;
  reg [16-1:0] _acc_0_x_source_generator_id;
  reg [32-1:0] _acc_0_x_source_offset;
  reg [33-1:0] _acc_0_x_source_size;
  reg [32-1:0] _acc_0_x_source_stride;
  reg [32-1:0] _acc_0_x_source_offset_buf;
  reg [33-1:0] _acc_0_x_source_size_buf;
  reg [32-1:0] _acc_0_x_source_stride_buf;
  reg [8-1:0] _acc_0_x_source_sel;
  reg [32-1:0] _acc_0_x_source_ram_raddr;
  reg _acc_0_x_source_ram_renable;
  wire [32-1:0] _acc_0_x_source_ram_rdata;
  reg _acc_0_x_source_fifo_deq;
  wire [32-1:0] _acc_0_x_source_fifo_rdata;
  reg [32-1:0] _acc_0_x_source_empty_data;
  reg _acc_0_rshift_idle;
  reg [33-1:0] _acc_0_rshift_source_count;
  reg [5-1:0] _acc_0_rshift_source_mode;
  reg [16-1:0] _acc_0_rshift_source_generator_id;
  reg [32-1:0] _acc_0_rshift_source_offset;
  reg [33-1:0] _acc_0_rshift_source_size;
  reg [32-1:0] _acc_0_rshift_source_stride;
  reg [32-1:0] _acc_0_rshift_source_offset_buf;
  reg [33-1:0] _acc_0_rshift_source_size_buf;
  reg [32-1:0] _acc_0_rshift_source_stride_buf;
  reg [8-1:0] _acc_0_rshift_source_sel;
  reg [32-1:0] _acc_0_rshift_source_ram_raddr;
  reg _acc_0_rshift_source_ram_renable;
  wire [32-1:0] _acc_0_rshift_source_ram_rdata;
  reg _acc_0_rshift_source_fifo_deq;
  wire [32-1:0] _acc_0_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_0_rshift_source_empty_data;
  reg [32-1:0] _acc_0_size_next_parameter_data;
  reg [33-1:0] _acc_0_sum_sink_count;
  reg [5-1:0] _acc_0_sum_sink_mode;
  reg [16-1:0] _acc_0_sum_sink_generator_id;
  reg [32-1:0] _acc_0_sum_sink_offset;
  reg [33-1:0] _acc_0_sum_sink_size;
  reg [32-1:0] _acc_0_sum_sink_stride;
  reg [32-1:0] _acc_0_sum_sink_offset_buf;
  reg [33-1:0] _acc_0_sum_sink_size_buf;
  reg [32-1:0] _acc_0_sum_sink_stride_buf;
  reg [8-1:0] _acc_0_sum_sink_sel;
  reg [32-1:0] _acc_0_sum_sink_waddr;
  reg _acc_0_sum_sink_wenable;
  reg [32-1:0] _acc_0_sum_sink_wdata;
  reg _acc_0_sum_sink_fifo_enq;
  reg [32-1:0] _acc_0_sum_sink_fifo_wdata;
  reg [32-1:0] _acc_0_sum_sink_immediate;
  reg [33-1:0] _acc_0_valid_sink_count;
  reg [5-1:0] _acc_0_valid_sink_mode;
  reg [16-1:0] _acc_0_valid_sink_generator_id;
  reg [32-1:0] _acc_0_valid_sink_offset;
  reg [33-1:0] _acc_0_valid_sink_size;
  reg [32-1:0] _acc_0_valid_sink_stride;
  reg [32-1:0] _acc_0_valid_sink_offset_buf;
  reg [33-1:0] _acc_0_valid_sink_size_buf;
  reg [32-1:0] _acc_0_valid_sink_stride_buf;
  reg [8-1:0] _acc_0_valid_sink_sel;
  reg [32-1:0] _acc_0_valid_sink_waddr;
  reg _acc_0_valid_sink_wenable;
  reg [1-1:0] _acc_0_valid_sink_wdata;
  reg _acc_0_valid_sink_fifo_enq;
  reg [1-1:0] _acc_0_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_0_valid_sink_immediate;
  reg _add_tree_1_stream_ivalid;
  wire _add_tree_1_stream_oready;
  wire _add_tree_1_stream_internal_oready;
  assign _add_tree_1_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_1_fsm;
  localparam _add_tree_1_fsm_init = 0;
  wire _add_tree_1_run_flag;
  assign _add_tree_1_run_flag = 0;
  reg _add_tree_1_source_start;
  wire _add_tree_1_source_stop;
  reg _add_tree_1_source_busy;
  wire _add_tree_1_sink_start;
  wire _add_tree_1_sink_stop;
  wire _add_tree_1_sink_busy;
  wire _add_tree_1_busy;
  reg _add_tree_1_busy_reg;
  wire _add_tree_1_is_root;
  reg _add_tree_1_var0_idle;
  reg [33-1:0] _add_tree_1_var0_source_count;
  reg [5-1:0] _add_tree_1_var0_source_mode;
  reg [16-1:0] _add_tree_1_var0_source_generator_id;
  reg [32-1:0] _add_tree_1_var0_source_offset;
  reg [33-1:0] _add_tree_1_var0_source_size;
  reg [32-1:0] _add_tree_1_var0_source_stride;
  reg [32-1:0] _add_tree_1_var0_source_offset_buf;
  reg [33-1:0] _add_tree_1_var0_source_size_buf;
  reg [32-1:0] _add_tree_1_var0_source_stride_buf;
  reg [8-1:0] _add_tree_1_var0_source_sel;
  reg [32-1:0] _add_tree_1_var0_source_ram_raddr;
  reg _add_tree_1_var0_source_ram_renable;
  wire [32-1:0] _add_tree_1_var0_source_ram_rdata;
  reg _add_tree_1_var0_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var0_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var0_source_empty_data;
  reg _add_tree_1_var1_idle;
  reg [33-1:0] _add_tree_1_var1_source_count;
  reg [5-1:0] _add_tree_1_var1_source_mode;
  reg [16-1:0] _add_tree_1_var1_source_generator_id;
  reg [32-1:0] _add_tree_1_var1_source_offset;
  reg [33-1:0] _add_tree_1_var1_source_size;
  reg [32-1:0] _add_tree_1_var1_source_stride;
  reg [32-1:0] _add_tree_1_var1_source_offset_buf;
  reg [33-1:0] _add_tree_1_var1_source_size_buf;
  reg [32-1:0] _add_tree_1_var1_source_stride_buf;
  reg [8-1:0] _add_tree_1_var1_source_sel;
  reg [32-1:0] _add_tree_1_var1_source_ram_raddr;
  reg _add_tree_1_var1_source_ram_renable;
  wire [32-1:0] _add_tree_1_var1_source_ram_rdata;
  reg _add_tree_1_var1_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var1_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var1_source_empty_data;
  reg _add_tree_1_var2_idle;
  reg [33-1:0] _add_tree_1_var2_source_count;
  reg [5-1:0] _add_tree_1_var2_source_mode;
  reg [16-1:0] _add_tree_1_var2_source_generator_id;
  reg [32-1:0] _add_tree_1_var2_source_offset;
  reg [33-1:0] _add_tree_1_var2_source_size;
  reg [32-1:0] _add_tree_1_var2_source_stride;
  reg [32-1:0] _add_tree_1_var2_source_offset_buf;
  reg [33-1:0] _add_tree_1_var2_source_size_buf;
  reg [32-1:0] _add_tree_1_var2_source_stride_buf;
  reg [8-1:0] _add_tree_1_var2_source_sel;
  reg [32-1:0] _add_tree_1_var2_source_ram_raddr;
  reg _add_tree_1_var2_source_ram_renable;
  wire [32-1:0] _add_tree_1_var2_source_ram_rdata;
  reg _add_tree_1_var2_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var2_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var2_source_empty_data;
  reg _add_tree_1_var3_idle;
  reg [33-1:0] _add_tree_1_var3_source_count;
  reg [5-1:0] _add_tree_1_var3_source_mode;
  reg [16-1:0] _add_tree_1_var3_source_generator_id;
  reg [32-1:0] _add_tree_1_var3_source_offset;
  reg [33-1:0] _add_tree_1_var3_source_size;
  reg [32-1:0] _add_tree_1_var3_source_stride;
  reg [32-1:0] _add_tree_1_var3_source_offset_buf;
  reg [33-1:0] _add_tree_1_var3_source_size_buf;
  reg [32-1:0] _add_tree_1_var3_source_stride_buf;
  reg [8-1:0] _add_tree_1_var3_source_sel;
  reg [32-1:0] _add_tree_1_var3_source_ram_raddr;
  reg _add_tree_1_var3_source_ram_renable;
  wire [32-1:0] _add_tree_1_var3_source_ram_rdata;
  reg _add_tree_1_var3_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var3_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var3_source_empty_data;
  reg _add_tree_1_var4_idle;
  reg [33-1:0] _add_tree_1_var4_source_count;
  reg [5-1:0] _add_tree_1_var4_source_mode;
  reg [16-1:0] _add_tree_1_var4_source_generator_id;
  reg [32-1:0] _add_tree_1_var4_source_offset;
  reg [33-1:0] _add_tree_1_var4_source_size;
  reg [32-1:0] _add_tree_1_var4_source_stride;
  reg [32-1:0] _add_tree_1_var4_source_offset_buf;
  reg [33-1:0] _add_tree_1_var4_source_size_buf;
  reg [32-1:0] _add_tree_1_var4_source_stride_buf;
  reg [8-1:0] _add_tree_1_var4_source_sel;
  reg [32-1:0] _add_tree_1_var4_source_ram_raddr;
  reg _add_tree_1_var4_source_ram_renable;
  wire [32-1:0] _add_tree_1_var4_source_ram_rdata;
  reg _add_tree_1_var4_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var4_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var4_source_empty_data;
  reg _add_tree_1_var5_idle;
  reg [33-1:0] _add_tree_1_var5_source_count;
  reg [5-1:0] _add_tree_1_var5_source_mode;
  reg [16-1:0] _add_tree_1_var5_source_generator_id;
  reg [32-1:0] _add_tree_1_var5_source_offset;
  reg [33-1:0] _add_tree_1_var5_source_size;
  reg [32-1:0] _add_tree_1_var5_source_stride;
  reg [32-1:0] _add_tree_1_var5_source_offset_buf;
  reg [33-1:0] _add_tree_1_var5_source_size_buf;
  reg [32-1:0] _add_tree_1_var5_source_stride_buf;
  reg [8-1:0] _add_tree_1_var5_source_sel;
  reg [32-1:0] _add_tree_1_var5_source_ram_raddr;
  reg _add_tree_1_var5_source_ram_renable;
  wire [32-1:0] _add_tree_1_var5_source_ram_rdata;
  reg _add_tree_1_var5_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var5_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var5_source_empty_data;
  reg _add_tree_1_var6_idle;
  reg [33-1:0] _add_tree_1_var6_source_count;
  reg [5-1:0] _add_tree_1_var6_source_mode;
  reg [16-1:0] _add_tree_1_var6_source_generator_id;
  reg [32-1:0] _add_tree_1_var6_source_offset;
  reg [33-1:0] _add_tree_1_var6_source_size;
  reg [32-1:0] _add_tree_1_var6_source_stride;
  reg [32-1:0] _add_tree_1_var6_source_offset_buf;
  reg [33-1:0] _add_tree_1_var6_source_size_buf;
  reg [32-1:0] _add_tree_1_var6_source_stride_buf;
  reg [8-1:0] _add_tree_1_var6_source_sel;
  reg [32-1:0] _add_tree_1_var6_source_ram_raddr;
  reg _add_tree_1_var6_source_ram_renable;
  wire [32-1:0] _add_tree_1_var6_source_ram_rdata;
  reg _add_tree_1_var6_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var6_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var6_source_empty_data;
  reg _add_tree_1_var7_idle;
  reg [33-1:0] _add_tree_1_var7_source_count;
  reg [5-1:0] _add_tree_1_var7_source_mode;
  reg [16-1:0] _add_tree_1_var7_source_generator_id;
  reg [32-1:0] _add_tree_1_var7_source_offset;
  reg [33-1:0] _add_tree_1_var7_source_size;
  reg [32-1:0] _add_tree_1_var7_source_stride;
  reg [32-1:0] _add_tree_1_var7_source_offset_buf;
  reg [33-1:0] _add_tree_1_var7_source_size_buf;
  reg [32-1:0] _add_tree_1_var7_source_stride_buf;
  reg [8-1:0] _add_tree_1_var7_source_sel;
  reg [32-1:0] _add_tree_1_var7_source_ram_raddr;
  reg _add_tree_1_var7_source_ram_renable;
  wire [32-1:0] _add_tree_1_var7_source_ram_rdata;
  reg _add_tree_1_var7_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var7_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var7_source_empty_data;
  reg _add_tree_1_var8_idle;
  reg [33-1:0] _add_tree_1_var8_source_count;
  reg [5-1:0] _add_tree_1_var8_source_mode;
  reg [16-1:0] _add_tree_1_var8_source_generator_id;
  reg [32-1:0] _add_tree_1_var8_source_offset;
  reg [33-1:0] _add_tree_1_var8_source_size;
  reg [32-1:0] _add_tree_1_var8_source_stride;
  reg [32-1:0] _add_tree_1_var8_source_offset_buf;
  reg [33-1:0] _add_tree_1_var8_source_size_buf;
  reg [32-1:0] _add_tree_1_var8_source_stride_buf;
  reg [8-1:0] _add_tree_1_var8_source_sel;
  reg [32-1:0] _add_tree_1_var8_source_ram_raddr;
  reg _add_tree_1_var8_source_ram_renable;
  wire [32-1:0] _add_tree_1_var8_source_ram_rdata;
  reg _add_tree_1_var8_source_fifo_deq;
  wire [32-1:0] _add_tree_1_var8_source_fifo_rdata;
  reg [32-1:0] _add_tree_1_var8_source_empty_data;
  reg [33-1:0] _add_tree_1_sum_sink_count;
  reg [5-1:0] _add_tree_1_sum_sink_mode;
  reg [16-1:0] _add_tree_1_sum_sink_generator_id;
  reg [32-1:0] _add_tree_1_sum_sink_offset;
  reg [33-1:0] _add_tree_1_sum_sink_size;
  reg [32-1:0] _add_tree_1_sum_sink_stride;
  reg [32-1:0] _add_tree_1_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_1_sum_sink_size_buf;
  reg [32-1:0] _add_tree_1_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_1_sum_sink_sel;
  reg [32-1:0] _add_tree_1_sum_sink_waddr;
  reg _add_tree_1_sum_sink_wenable;
  reg [32-1:0] _add_tree_1_sum_sink_wdata;
  reg _add_tree_1_sum_sink_fifo_enq;
  reg [32-1:0] _add_tree_1_sum_sink_fifo_wdata;
  reg [32-1:0] _add_tree_1_sum_sink_immediate;
  reg _mul_rshift_round_clip_2_stream_ivalid;
  wire _mul_rshift_round_clip_2_stream_oready;
  wire _mul_rshift_round_clip_2_stream_internal_oready;
  assign _mul_rshift_round_clip_2_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_2_fsm;
  localparam _mul_rshift_round_clip_2_fsm_init = 0;
  wire _mul_rshift_round_clip_2_run_flag;
  assign _mul_rshift_round_clip_2_run_flag = 0;
  reg _mul_rshift_round_clip_2_source_start;
  wire _mul_rshift_round_clip_2_source_stop;
  reg _mul_rshift_round_clip_2_source_busy;
  wire _mul_rshift_round_clip_2_sink_start;
  wire _mul_rshift_round_clip_2_sink_stop;
  wire _mul_rshift_round_clip_2_sink_busy;
  wire _mul_rshift_round_clip_2_busy;
  reg _mul_rshift_round_clip_2_busy_reg;
  wire _mul_rshift_round_clip_2_is_root;
  reg _mul_rshift_round_clip_2_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_2_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_2_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_2_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_2_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_2_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_2_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_2_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_2_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_2_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_2_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_2_x_source_ram_raddr;
  reg _mul_rshift_round_clip_2_x_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_2_x_source_ram_rdata;
  reg _mul_rshift_round_clip_2_x_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_2_x_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_2_x_source_empty_data;
  reg _mul_rshift_round_clip_2_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_2_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_2_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_2_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_2_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_2_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_2_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_2_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_2_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_2_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_2_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_2_y_source_ram_raddr;
  reg _mul_rshift_round_clip_2_y_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_2_y_source_ram_rdata;
  reg _mul_rshift_round_clip_2_y_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_2_y_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_2_y_source_empty_data;
  reg _mul_rshift_round_clip_2_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_2_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_2_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_2_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_2_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_2_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_2_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_2_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_2_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_2_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_2_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_2_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_2_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_2_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_2_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_2_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_2_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_2_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_2_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_2_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_2_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_2_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_2_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_waddr;
  reg _mul_rshift_round_clip_2_z_sink_wenable;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_wdata;
  reg _mul_rshift_round_clip_2_z_sink_fifo_enq;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_fifo_wdata;
  reg [32-1:0] _mul_rshift_round_clip_2_z_sink_immediate;
  reg _mul_3_stream_ivalid;
  wire _mul_3_stream_oready;
  wire _mul_3_stream_internal_oready;
  assign _mul_3_stream_internal_oready = 1;
  reg [32-1:0] _mul_3_fsm;
  localparam _mul_3_fsm_init = 0;
  wire _mul_3_run_flag;
  assign _mul_3_run_flag = 0;
  reg _mul_3_source_start;
  wire _mul_3_source_stop;
  reg _mul_3_source_busy;
  wire _mul_3_sink_start;
  wire _mul_3_sink_stop;
  wire _mul_3_sink_busy;
  wire _mul_3_busy;
  reg _mul_3_busy_reg;
  wire _mul_3_is_root;
  reg _mul_3_x_idle;
  reg [33-1:0] _mul_3_x_source_count;
  reg [5-1:0] _mul_3_x_source_mode;
  reg [16-1:0] _mul_3_x_source_generator_id;
  reg [32-1:0] _mul_3_x_source_offset;
  reg [33-1:0] _mul_3_x_source_size;
  reg [32-1:0] _mul_3_x_source_stride;
  reg [32-1:0] _mul_3_x_source_offset_buf;
  reg [33-1:0] _mul_3_x_source_size_buf;
  reg [32-1:0] _mul_3_x_source_stride_buf;
  reg [8-1:0] _mul_3_x_source_sel;
  reg [32-1:0] _mul_3_x_source_ram_raddr;
  reg _mul_3_x_source_ram_renable;
  wire [32-1:0] _mul_3_x_source_ram_rdata;
  reg _mul_3_x_source_fifo_deq;
  wire [32-1:0] _mul_3_x_source_fifo_rdata;
  reg [32-1:0] _mul_3_x_source_empty_data;
  reg _mul_3_y_idle;
  reg [33-1:0] _mul_3_y_source_count;
  reg [5-1:0] _mul_3_y_source_mode;
  reg [16-1:0] _mul_3_y_source_generator_id;
  reg [32-1:0] _mul_3_y_source_offset;
  reg [33-1:0] _mul_3_y_source_size;
  reg [32-1:0] _mul_3_y_source_stride;
  reg [32-1:0] _mul_3_y_source_offset_buf;
  reg [33-1:0] _mul_3_y_source_size_buf;
  reg [32-1:0] _mul_3_y_source_stride_buf;
  reg [8-1:0] _mul_3_y_source_sel;
  reg [32-1:0] _mul_3_y_source_ram_raddr;
  reg _mul_3_y_source_ram_renable;
  wire [32-1:0] _mul_3_y_source_ram_rdata;
  reg _mul_3_y_source_fifo_deq;
  wire [32-1:0] _mul_3_y_source_fifo_rdata;
  reg [32-1:0] _mul_3_y_source_empty_data;
  reg _mul_3_rshift_idle;
  reg [33-1:0] _mul_3_rshift_source_count;
  reg [5-1:0] _mul_3_rshift_source_mode;
  reg [16-1:0] _mul_3_rshift_source_generator_id;
  reg [32-1:0] _mul_3_rshift_source_offset;
  reg [33-1:0] _mul_3_rshift_source_size;
  reg [32-1:0] _mul_3_rshift_source_stride;
  reg [32-1:0] _mul_3_rshift_source_offset_buf;
  reg [33-1:0] _mul_3_rshift_source_size_buf;
  reg [32-1:0] _mul_3_rshift_source_stride_buf;
  reg [8-1:0] _mul_3_rshift_source_sel;
  reg [32-1:0] _mul_3_rshift_source_ram_raddr;
  reg _mul_3_rshift_source_ram_renable;
  wire [32-1:0] _mul_3_rshift_source_ram_rdata;
  reg _mul_3_rshift_source_fifo_deq;
  wire [32-1:0] _mul_3_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_3_rshift_source_empty_data;
  reg [33-1:0] _mul_3_z_sink_count;
  reg [5-1:0] _mul_3_z_sink_mode;
  reg [16-1:0] _mul_3_z_sink_generator_id;
  reg [32-1:0] _mul_3_z_sink_offset;
  reg [33-1:0] _mul_3_z_sink_size;
  reg [32-1:0] _mul_3_z_sink_stride;
  reg [32-1:0] _mul_3_z_sink_offset_buf;
  reg [33-1:0] _mul_3_z_sink_size_buf;
  reg [32-1:0] _mul_3_z_sink_stride_buf;
  reg [8-1:0] _mul_3_z_sink_sel;
  reg [32-1:0] _mul_3_z_sink_waddr;
  reg _mul_3_z_sink_wenable;
  reg [32-1:0] _mul_3_z_sink_wdata;
  reg _mul_3_z_sink_fifo_enq;
  reg [32-1:0] _mul_3_z_sink_fifo_wdata;
  reg [32-1:0] _mul_3_z_sink_immediate;
  reg _mul_4_stream_ivalid;
  wire _mul_4_stream_oready;
  wire _mul_4_stream_internal_oready;
  assign _mul_4_stream_internal_oready = 1;
  reg [32-1:0] _mul_4_fsm;
  localparam _mul_4_fsm_init = 0;
  wire _mul_4_run_flag;
  assign _mul_4_run_flag = 0;
  reg _mul_4_source_start;
  wire _mul_4_source_stop;
  reg _mul_4_source_busy;
  wire _mul_4_sink_start;
  wire _mul_4_sink_stop;
  wire _mul_4_sink_busy;
  wire _mul_4_busy;
  reg _mul_4_busy_reg;
  wire _mul_4_is_root;
  reg _mul_4_x_idle;
  reg [33-1:0] _mul_4_x_source_count;
  reg [5-1:0] _mul_4_x_source_mode;
  reg [16-1:0] _mul_4_x_source_generator_id;
  reg [32-1:0] _mul_4_x_source_offset;
  reg [33-1:0] _mul_4_x_source_size;
  reg [32-1:0] _mul_4_x_source_stride;
  reg [32-1:0] _mul_4_x_source_offset_buf;
  reg [33-1:0] _mul_4_x_source_size_buf;
  reg [32-1:0] _mul_4_x_source_stride_buf;
  reg [8-1:0] _mul_4_x_source_sel;
  reg [32-1:0] _mul_4_x_source_ram_raddr;
  reg _mul_4_x_source_ram_renable;
  wire [32-1:0] _mul_4_x_source_ram_rdata;
  reg _mul_4_x_source_fifo_deq;
  wire [32-1:0] _mul_4_x_source_fifo_rdata;
  reg [32-1:0] _mul_4_x_source_empty_data;
  reg _mul_4_y_idle;
  reg [33-1:0] _mul_4_y_source_count;
  reg [5-1:0] _mul_4_y_source_mode;
  reg [16-1:0] _mul_4_y_source_generator_id;
  reg [32-1:0] _mul_4_y_source_offset;
  reg [33-1:0] _mul_4_y_source_size;
  reg [32-1:0] _mul_4_y_source_stride;
  reg [32-1:0] _mul_4_y_source_offset_buf;
  reg [33-1:0] _mul_4_y_source_size_buf;
  reg [32-1:0] _mul_4_y_source_stride_buf;
  reg [8-1:0] _mul_4_y_source_sel;
  reg [32-1:0] _mul_4_y_source_ram_raddr;
  reg _mul_4_y_source_ram_renable;
  wire [32-1:0] _mul_4_y_source_ram_rdata;
  reg _mul_4_y_source_fifo_deq;
  wire [32-1:0] _mul_4_y_source_fifo_rdata;
  reg [32-1:0] _mul_4_y_source_empty_data;
  reg _mul_4_rshift_idle;
  reg [33-1:0] _mul_4_rshift_source_count;
  reg [5-1:0] _mul_4_rshift_source_mode;
  reg [16-1:0] _mul_4_rshift_source_generator_id;
  reg [32-1:0] _mul_4_rshift_source_offset;
  reg [33-1:0] _mul_4_rshift_source_size;
  reg [32-1:0] _mul_4_rshift_source_stride;
  reg [32-1:0] _mul_4_rshift_source_offset_buf;
  reg [33-1:0] _mul_4_rshift_source_size_buf;
  reg [32-1:0] _mul_4_rshift_source_stride_buf;
  reg [8-1:0] _mul_4_rshift_source_sel;
  reg [32-1:0] _mul_4_rshift_source_ram_raddr;
  reg _mul_4_rshift_source_ram_renable;
  wire [32-1:0] _mul_4_rshift_source_ram_rdata;
  reg _mul_4_rshift_source_fifo_deq;
  wire [32-1:0] _mul_4_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_4_rshift_source_empty_data;
  reg [33-1:0] _mul_4_z_sink_count;
  reg [5-1:0] _mul_4_z_sink_mode;
  reg [16-1:0] _mul_4_z_sink_generator_id;
  reg [32-1:0] _mul_4_z_sink_offset;
  reg [33-1:0] _mul_4_z_sink_size;
  reg [32-1:0] _mul_4_z_sink_stride;
  reg [32-1:0] _mul_4_z_sink_offset_buf;
  reg [33-1:0] _mul_4_z_sink_size_buf;
  reg [32-1:0] _mul_4_z_sink_stride_buf;
  reg [8-1:0] _mul_4_z_sink_sel;
  reg [32-1:0] _mul_4_z_sink_waddr;
  reg _mul_4_z_sink_wenable;
  reg [32-1:0] _mul_4_z_sink_wdata;
  reg _mul_4_z_sink_fifo_enq;
  reg [32-1:0] _mul_4_z_sink_fifo_wdata;
  reg [32-1:0] _mul_4_z_sink_immediate;
  reg _mul_5_stream_ivalid;
  wire _mul_5_stream_oready;
  wire _mul_5_stream_internal_oready;
  assign _mul_5_stream_internal_oready = 1;
  reg [32-1:0] _mul_5_fsm;
  localparam _mul_5_fsm_init = 0;
  wire _mul_5_run_flag;
  assign _mul_5_run_flag = 0;
  reg _mul_5_source_start;
  wire _mul_5_source_stop;
  reg _mul_5_source_busy;
  wire _mul_5_sink_start;
  wire _mul_5_sink_stop;
  wire _mul_5_sink_busy;
  wire _mul_5_busy;
  reg _mul_5_busy_reg;
  wire _mul_5_is_root;
  reg _mul_5_x_idle;
  reg [33-1:0] _mul_5_x_source_count;
  reg [5-1:0] _mul_5_x_source_mode;
  reg [16-1:0] _mul_5_x_source_generator_id;
  reg [32-1:0] _mul_5_x_source_offset;
  reg [33-1:0] _mul_5_x_source_size;
  reg [32-1:0] _mul_5_x_source_stride;
  reg [32-1:0] _mul_5_x_source_offset_buf;
  reg [33-1:0] _mul_5_x_source_size_buf;
  reg [32-1:0] _mul_5_x_source_stride_buf;
  reg [8-1:0] _mul_5_x_source_sel;
  reg [32-1:0] _mul_5_x_source_ram_raddr;
  reg _mul_5_x_source_ram_renable;
  wire [32-1:0] _mul_5_x_source_ram_rdata;
  reg _mul_5_x_source_fifo_deq;
  wire [32-1:0] _mul_5_x_source_fifo_rdata;
  reg [32-1:0] _mul_5_x_source_empty_data;
  reg _mul_5_y_idle;
  reg [33-1:0] _mul_5_y_source_count;
  reg [5-1:0] _mul_5_y_source_mode;
  reg [16-1:0] _mul_5_y_source_generator_id;
  reg [32-1:0] _mul_5_y_source_offset;
  reg [33-1:0] _mul_5_y_source_size;
  reg [32-1:0] _mul_5_y_source_stride;
  reg [32-1:0] _mul_5_y_source_offset_buf;
  reg [33-1:0] _mul_5_y_source_size_buf;
  reg [32-1:0] _mul_5_y_source_stride_buf;
  reg [8-1:0] _mul_5_y_source_sel;
  reg [32-1:0] _mul_5_y_source_ram_raddr;
  reg _mul_5_y_source_ram_renable;
  wire [32-1:0] _mul_5_y_source_ram_rdata;
  reg _mul_5_y_source_fifo_deq;
  wire [32-1:0] _mul_5_y_source_fifo_rdata;
  reg [32-1:0] _mul_5_y_source_empty_data;
  reg _mul_5_rshift_idle;
  reg [33-1:0] _mul_5_rshift_source_count;
  reg [5-1:0] _mul_5_rshift_source_mode;
  reg [16-1:0] _mul_5_rshift_source_generator_id;
  reg [32-1:0] _mul_5_rshift_source_offset;
  reg [33-1:0] _mul_5_rshift_source_size;
  reg [32-1:0] _mul_5_rshift_source_stride;
  reg [32-1:0] _mul_5_rshift_source_offset_buf;
  reg [33-1:0] _mul_5_rshift_source_size_buf;
  reg [32-1:0] _mul_5_rshift_source_stride_buf;
  reg [8-1:0] _mul_5_rshift_source_sel;
  reg [32-1:0] _mul_5_rshift_source_ram_raddr;
  reg _mul_5_rshift_source_ram_renable;
  wire [32-1:0] _mul_5_rshift_source_ram_rdata;
  reg _mul_5_rshift_source_fifo_deq;
  wire [32-1:0] _mul_5_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_5_rshift_source_empty_data;
  reg [33-1:0] _mul_5_z_sink_count;
  reg [5-1:0] _mul_5_z_sink_mode;
  reg [16-1:0] _mul_5_z_sink_generator_id;
  reg [32-1:0] _mul_5_z_sink_offset;
  reg [33-1:0] _mul_5_z_sink_size;
  reg [32-1:0] _mul_5_z_sink_stride;
  reg [32-1:0] _mul_5_z_sink_offset_buf;
  reg [33-1:0] _mul_5_z_sink_size_buf;
  reg [32-1:0] _mul_5_z_sink_stride_buf;
  reg [8-1:0] _mul_5_z_sink_sel;
  reg [32-1:0] _mul_5_z_sink_waddr;
  reg _mul_5_z_sink_wenable;
  reg [32-1:0] _mul_5_z_sink_wdata;
  reg _mul_5_z_sink_fifo_enq;
  reg [32-1:0] _mul_5_z_sink_fifo_wdata;
  reg [32-1:0] _mul_5_z_sink_immediate;
  reg _mul_6_stream_ivalid;
  wire _mul_6_stream_oready;
  wire _mul_6_stream_internal_oready;
  assign _mul_6_stream_internal_oready = 1;
  reg [32-1:0] _mul_6_fsm;
  localparam _mul_6_fsm_init = 0;
  wire _mul_6_run_flag;
  assign _mul_6_run_flag = 0;
  reg _mul_6_source_start;
  wire _mul_6_source_stop;
  reg _mul_6_source_busy;
  wire _mul_6_sink_start;
  wire _mul_6_sink_stop;
  wire _mul_6_sink_busy;
  wire _mul_6_busy;
  reg _mul_6_busy_reg;
  wire _mul_6_is_root;
  reg _mul_6_x_idle;
  reg [33-1:0] _mul_6_x_source_count;
  reg [5-1:0] _mul_6_x_source_mode;
  reg [16-1:0] _mul_6_x_source_generator_id;
  reg [32-1:0] _mul_6_x_source_offset;
  reg [33-1:0] _mul_6_x_source_size;
  reg [32-1:0] _mul_6_x_source_stride;
  reg [32-1:0] _mul_6_x_source_offset_buf;
  reg [33-1:0] _mul_6_x_source_size_buf;
  reg [32-1:0] _mul_6_x_source_stride_buf;
  reg [8-1:0] _mul_6_x_source_sel;
  reg [32-1:0] _mul_6_x_source_ram_raddr;
  reg _mul_6_x_source_ram_renable;
  wire [32-1:0] _mul_6_x_source_ram_rdata;
  reg _mul_6_x_source_fifo_deq;
  wire [32-1:0] _mul_6_x_source_fifo_rdata;
  reg [32-1:0] _mul_6_x_source_empty_data;
  reg _mul_6_y_idle;
  reg [33-1:0] _mul_6_y_source_count;
  reg [5-1:0] _mul_6_y_source_mode;
  reg [16-1:0] _mul_6_y_source_generator_id;
  reg [32-1:0] _mul_6_y_source_offset;
  reg [33-1:0] _mul_6_y_source_size;
  reg [32-1:0] _mul_6_y_source_stride;
  reg [32-1:0] _mul_6_y_source_offset_buf;
  reg [33-1:0] _mul_6_y_source_size_buf;
  reg [32-1:0] _mul_6_y_source_stride_buf;
  reg [8-1:0] _mul_6_y_source_sel;
  reg [32-1:0] _mul_6_y_source_ram_raddr;
  reg _mul_6_y_source_ram_renable;
  wire [32-1:0] _mul_6_y_source_ram_rdata;
  reg _mul_6_y_source_fifo_deq;
  wire [32-1:0] _mul_6_y_source_fifo_rdata;
  reg [32-1:0] _mul_6_y_source_empty_data;
  reg _mul_6_rshift_idle;
  reg [33-1:0] _mul_6_rshift_source_count;
  reg [5-1:0] _mul_6_rshift_source_mode;
  reg [16-1:0] _mul_6_rshift_source_generator_id;
  reg [32-1:0] _mul_6_rshift_source_offset;
  reg [33-1:0] _mul_6_rshift_source_size;
  reg [32-1:0] _mul_6_rshift_source_stride;
  reg [32-1:0] _mul_6_rshift_source_offset_buf;
  reg [33-1:0] _mul_6_rshift_source_size_buf;
  reg [32-1:0] _mul_6_rshift_source_stride_buf;
  reg [8-1:0] _mul_6_rshift_source_sel;
  reg [32-1:0] _mul_6_rshift_source_ram_raddr;
  reg _mul_6_rshift_source_ram_renable;
  wire [32-1:0] _mul_6_rshift_source_ram_rdata;
  reg _mul_6_rshift_source_fifo_deq;
  wire [32-1:0] _mul_6_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_6_rshift_source_empty_data;
  reg [33-1:0] _mul_6_z_sink_count;
  reg [5-1:0] _mul_6_z_sink_mode;
  reg [16-1:0] _mul_6_z_sink_generator_id;
  reg [32-1:0] _mul_6_z_sink_offset;
  reg [33-1:0] _mul_6_z_sink_size;
  reg [32-1:0] _mul_6_z_sink_stride;
  reg [32-1:0] _mul_6_z_sink_offset_buf;
  reg [33-1:0] _mul_6_z_sink_size_buf;
  reg [32-1:0] _mul_6_z_sink_stride_buf;
  reg [8-1:0] _mul_6_z_sink_sel;
  reg [32-1:0] _mul_6_z_sink_waddr;
  reg _mul_6_z_sink_wenable;
  reg [32-1:0] _mul_6_z_sink_wdata;
  reg _mul_6_z_sink_fifo_enq;
  reg [32-1:0] _mul_6_z_sink_fifo_wdata;
  reg [32-1:0] _mul_6_z_sink_immediate;
  reg _mul_7_stream_ivalid;
  wire _mul_7_stream_oready;
  wire _mul_7_stream_internal_oready;
  assign _mul_7_stream_internal_oready = 1;
  reg [32-1:0] _mul_7_fsm;
  localparam _mul_7_fsm_init = 0;
  wire _mul_7_run_flag;
  assign _mul_7_run_flag = 0;
  reg _mul_7_source_start;
  wire _mul_7_source_stop;
  reg _mul_7_source_busy;
  wire _mul_7_sink_start;
  wire _mul_7_sink_stop;
  wire _mul_7_sink_busy;
  wire _mul_7_busy;
  reg _mul_7_busy_reg;
  wire _mul_7_is_root;
  reg _mul_7_x_idle;
  reg [33-1:0] _mul_7_x_source_count;
  reg [5-1:0] _mul_7_x_source_mode;
  reg [16-1:0] _mul_7_x_source_generator_id;
  reg [32-1:0] _mul_7_x_source_offset;
  reg [33-1:0] _mul_7_x_source_size;
  reg [32-1:0] _mul_7_x_source_stride;
  reg [32-1:0] _mul_7_x_source_offset_buf;
  reg [33-1:0] _mul_7_x_source_size_buf;
  reg [32-1:0] _mul_7_x_source_stride_buf;
  reg [8-1:0] _mul_7_x_source_sel;
  reg [32-1:0] _mul_7_x_source_ram_raddr;
  reg _mul_7_x_source_ram_renable;
  wire [32-1:0] _mul_7_x_source_ram_rdata;
  reg _mul_7_x_source_fifo_deq;
  wire [32-1:0] _mul_7_x_source_fifo_rdata;
  reg [32-1:0] _mul_7_x_source_empty_data;
  reg _mul_7_y_idle;
  reg [33-1:0] _mul_7_y_source_count;
  reg [5-1:0] _mul_7_y_source_mode;
  reg [16-1:0] _mul_7_y_source_generator_id;
  reg [32-1:0] _mul_7_y_source_offset;
  reg [33-1:0] _mul_7_y_source_size;
  reg [32-1:0] _mul_7_y_source_stride;
  reg [32-1:0] _mul_7_y_source_offset_buf;
  reg [33-1:0] _mul_7_y_source_size_buf;
  reg [32-1:0] _mul_7_y_source_stride_buf;
  reg [8-1:0] _mul_7_y_source_sel;
  reg [32-1:0] _mul_7_y_source_ram_raddr;
  reg _mul_7_y_source_ram_renable;
  wire [32-1:0] _mul_7_y_source_ram_rdata;
  reg _mul_7_y_source_fifo_deq;
  wire [32-1:0] _mul_7_y_source_fifo_rdata;
  reg [32-1:0] _mul_7_y_source_empty_data;
  reg _mul_7_rshift_idle;
  reg [33-1:0] _mul_7_rshift_source_count;
  reg [5-1:0] _mul_7_rshift_source_mode;
  reg [16-1:0] _mul_7_rshift_source_generator_id;
  reg [32-1:0] _mul_7_rshift_source_offset;
  reg [33-1:0] _mul_7_rshift_source_size;
  reg [32-1:0] _mul_7_rshift_source_stride;
  reg [32-1:0] _mul_7_rshift_source_offset_buf;
  reg [33-1:0] _mul_7_rshift_source_size_buf;
  reg [32-1:0] _mul_7_rshift_source_stride_buf;
  reg [8-1:0] _mul_7_rshift_source_sel;
  reg [32-1:0] _mul_7_rshift_source_ram_raddr;
  reg _mul_7_rshift_source_ram_renable;
  wire [32-1:0] _mul_7_rshift_source_ram_rdata;
  reg _mul_7_rshift_source_fifo_deq;
  wire [32-1:0] _mul_7_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_7_rshift_source_empty_data;
  reg [33-1:0] _mul_7_z_sink_count;
  reg [5-1:0] _mul_7_z_sink_mode;
  reg [16-1:0] _mul_7_z_sink_generator_id;
  reg [32-1:0] _mul_7_z_sink_offset;
  reg [33-1:0] _mul_7_z_sink_size;
  reg [32-1:0] _mul_7_z_sink_stride;
  reg [32-1:0] _mul_7_z_sink_offset_buf;
  reg [33-1:0] _mul_7_z_sink_size_buf;
  reg [32-1:0] _mul_7_z_sink_stride_buf;
  reg [8-1:0] _mul_7_z_sink_sel;
  reg [32-1:0] _mul_7_z_sink_waddr;
  reg _mul_7_z_sink_wenable;
  reg [32-1:0] _mul_7_z_sink_wdata;
  reg _mul_7_z_sink_fifo_enq;
  reg [32-1:0] _mul_7_z_sink_fifo_wdata;
  reg [32-1:0] _mul_7_z_sink_immediate;
  reg _mul_8_stream_ivalid;
  wire _mul_8_stream_oready;
  wire _mul_8_stream_internal_oready;
  assign _mul_8_stream_internal_oready = 1;
  reg [32-1:0] _mul_8_fsm;
  localparam _mul_8_fsm_init = 0;
  wire _mul_8_run_flag;
  assign _mul_8_run_flag = 0;
  reg _mul_8_source_start;
  wire _mul_8_source_stop;
  reg _mul_8_source_busy;
  wire _mul_8_sink_start;
  wire _mul_8_sink_stop;
  wire _mul_8_sink_busy;
  wire _mul_8_busy;
  reg _mul_8_busy_reg;
  wire _mul_8_is_root;
  reg _mul_8_x_idle;
  reg [33-1:0] _mul_8_x_source_count;
  reg [5-1:0] _mul_8_x_source_mode;
  reg [16-1:0] _mul_8_x_source_generator_id;
  reg [32-1:0] _mul_8_x_source_offset;
  reg [33-1:0] _mul_8_x_source_size;
  reg [32-1:0] _mul_8_x_source_stride;
  reg [32-1:0] _mul_8_x_source_offset_buf;
  reg [33-1:0] _mul_8_x_source_size_buf;
  reg [32-1:0] _mul_8_x_source_stride_buf;
  reg [8-1:0] _mul_8_x_source_sel;
  reg [32-1:0] _mul_8_x_source_ram_raddr;
  reg _mul_8_x_source_ram_renable;
  wire [32-1:0] _mul_8_x_source_ram_rdata;
  reg _mul_8_x_source_fifo_deq;
  wire [32-1:0] _mul_8_x_source_fifo_rdata;
  reg [32-1:0] _mul_8_x_source_empty_data;
  reg _mul_8_y_idle;
  reg [33-1:0] _mul_8_y_source_count;
  reg [5-1:0] _mul_8_y_source_mode;
  reg [16-1:0] _mul_8_y_source_generator_id;
  reg [32-1:0] _mul_8_y_source_offset;
  reg [33-1:0] _mul_8_y_source_size;
  reg [32-1:0] _mul_8_y_source_stride;
  reg [32-1:0] _mul_8_y_source_offset_buf;
  reg [33-1:0] _mul_8_y_source_size_buf;
  reg [32-1:0] _mul_8_y_source_stride_buf;
  reg [8-1:0] _mul_8_y_source_sel;
  reg [32-1:0] _mul_8_y_source_ram_raddr;
  reg _mul_8_y_source_ram_renable;
  wire [32-1:0] _mul_8_y_source_ram_rdata;
  reg _mul_8_y_source_fifo_deq;
  wire [32-1:0] _mul_8_y_source_fifo_rdata;
  reg [32-1:0] _mul_8_y_source_empty_data;
  reg _mul_8_rshift_idle;
  reg [33-1:0] _mul_8_rshift_source_count;
  reg [5-1:0] _mul_8_rshift_source_mode;
  reg [16-1:0] _mul_8_rshift_source_generator_id;
  reg [32-1:0] _mul_8_rshift_source_offset;
  reg [33-1:0] _mul_8_rshift_source_size;
  reg [32-1:0] _mul_8_rshift_source_stride;
  reg [32-1:0] _mul_8_rshift_source_offset_buf;
  reg [33-1:0] _mul_8_rshift_source_size_buf;
  reg [32-1:0] _mul_8_rshift_source_stride_buf;
  reg [8-1:0] _mul_8_rshift_source_sel;
  reg [32-1:0] _mul_8_rshift_source_ram_raddr;
  reg _mul_8_rshift_source_ram_renable;
  wire [32-1:0] _mul_8_rshift_source_ram_rdata;
  reg _mul_8_rshift_source_fifo_deq;
  wire [32-1:0] _mul_8_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_8_rshift_source_empty_data;
  reg [33-1:0] _mul_8_z_sink_count;
  reg [5-1:0] _mul_8_z_sink_mode;
  reg [16-1:0] _mul_8_z_sink_generator_id;
  reg [32-1:0] _mul_8_z_sink_offset;
  reg [33-1:0] _mul_8_z_sink_size;
  reg [32-1:0] _mul_8_z_sink_stride;
  reg [32-1:0] _mul_8_z_sink_offset_buf;
  reg [33-1:0] _mul_8_z_sink_size_buf;
  reg [32-1:0] _mul_8_z_sink_stride_buf;
  reg [8-1:0] _mul_8_z_sink_sel;
  reg [32-1:0] _mul_8_z_sink_waddr;
  reg _mul_8_z_sink_wenable;
  reg [32-1:0] _mul_8_z_sink_wdata;
  reg _mul_8_z_sink_fifo_enq;
  reg [32-1:0] _mul_8_z_sink_fifo_wdata;
  reg [32-1:0] _mul_8_z_sink_immediate;
  reg _mul_9_stream_ivalid;
  wire _mul_9_stream_oready;
  wire _mul_9_stream_internal_oready;
  assign _mul_9_stream_internal_oready = 1;
  reg [32-1:0] _mul_9_fsm;
  localparam _mul_9_fsm_init = 0;
  wire _mul_9_run_flag;
  assign _mul_9_run_flag = 0;
  reg _mul_9_source_start;
  wire _mul_9_source_stop;
  reg _mul_9_source_busy;
  wire _mul_9_sink_start;
  wire _mul_9_sink_stop;
  wire _mul_9_sink_busy;
  wire _mul_9_busy;
  reg _mul_9_busy_reg;
  wire _mul_9_is_root;
  reg _mul_9_x_idle;
  reg [33-1:0] _mul_9_x_source_count;
  reg [5-1:0] _mul_9_x_source_mode;
  reg [16-1:0] _mul_9_x_source_generator_id;
  reg [32-1:0] _mul_9_x_source_offset;
  reg [33-1:0] _mul_9_x_source_size;
  reg [32-1:0] _mul_9_x_source_stride;
  reg [32-1:0] _mul_9_x_source_offset_buf;
  reg [33-1:0] _mul_9_x_source_size_buf;
  reg [32-1:0] _mul_9_x_source_stride_buf;
  reg [8-1:0] _mul_9_x_source_sel;
  reg [32-1:0] _mul_9_x_source_ram_raddr;
  reg _mul_9_x_source_ram_renable;
  wire [32-1:0] _mul_9_x_source_ram_rdata;
  reg _mul_9_x_source_fifo_deq;
  wire [32-1:0] _mul_9_x_source_fifo_rdata;
  reg [32-1:0] _mul_9_x_source_empty_data;
  reg _mul_9_y_idle;
  reg [33-1:0] _mul_9_y_source_count;
  reg [5-1:0] _mul_9_y_source_mode;
  reg [16-1:0] _mul_9_y_source_generator_id;
  reg [32-1:0] _mul_9_y_source_offset;
  reg [33-1:0] _mul_9_y_source_size;
  reg [32-1:0] _mul_9_y_source_stride;
  reg [32-1:0] _mul_9_y_source_offset_buf;
  reg [33-1:0] _mul_9_y_source_size_buf;
  reg [32-1:0] _mul_9_y_source_stride_buf;
  reg [8-1:0] _mul_9_y_source_sel;
  reg [32-1:0] _mul_9_y_source_ram_raddr;
  reg _mul_9_y_source_ram_renable;
  wire [32-1:0] _mul_9_y_source_ram_rdata;
  reg _mul_9_y_source_fifo_deq;
  wire [32-1:0] _mul_9_y_source_fifo_rdata;
  reg [32-1:0] _mul_9_y_source_empty_data;
  reg _mul_9_rshift_idle;
  reg [33-1:0] _mul_9_rshift_source_count;
  reg [5-1:0] _mul_9_rshift_source_mode;
  reg [16-1:0] _mul_9_rshift_source_generator_id;
  reg [32-1:0] _mul_9_rshift_source_offset;
  reg [33-1:0] _mul_9_rshift_source_size;
  reg [32-1:0] _mul_9_rshift_source_stride;
  reg [32-1:0] _mul_9_rshift_source_offset_buf;
  reg [33-1:0] _mul_9_rshift_source_size_buf;
  reg [32-1:0] _mul_9_rshift_source_stride_buf;
  reg [8-1:0] _mul_9_rshift_source_sel;
  reg [32-1:0] _mul_9_rshift_source_ram_raddr;
  reg _mul_9_rshift_source_ram_renable;
  wire [32-1:0] _mul_9_rshift_source_ram_rdata;
  reg _mul_9_rshift_source_fifo_deq;
  wire [32-1:0] _mul_9_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_9_rshift_source_empty_data;
  reg [33-1:0] _mul_9_z_sink_count;
  reg [5-1:0] _mul_9_z_sink_mode;
  reg [16-1:0] _mul_9_z_sink_generator_id;
  reg [32-1:0] _mul_9_z_sink_offset;
  reg [33-1:0] _mul_9_z_sink_size;
  reg [32-1:0] _mul_9_z_sink_stride;
  reg [32-1:0] _mul_9_z_sink_offset_buf;
  reg [33-1:0] _mul_9_z_sink_size_buf;
  reg [32-1:0] _mul_9_z_sink_stride_buf;
  reg [8-1:0] _mul_9_z_sink_sel;
  reg [32-1:0] _mul_9_z_sink_waddr;
  reg _mul_9_z_sink_wenable;
  reg [32-1:0] _mul_9_z_sink_wdata;
  reg _mul_9_z_sink_fifo_enq;
  reg [32-1:0] _mul_9_z_sink_fifo_wdata;
  reg [32-1:0] _mul_9_z_sink_immediate;
  reg _mul_10_stream_ivalid;
  wire _mul_10_stream_oready;
  wire _mul_10_stream_internal_oready;
  assign _mul_10_stream_internal_oready = 1;
  reg [32-1:0] _mul_10_fsm;
  localparam _mul_10_fsm_init = 0;
  wire _mul_10_run_flag;
  assign _mul_10_run_flag = 0;
  reg _mul_10_source_start;
  wire _mul_10_source_stop;
  reg _mul_10_source_busy;
  wire _mul_10_sink_start;
  wire _mul_10_sink_stop;
  wire _mul_10_sink_busy;
  wire _mul_10_busy;
  reg _mul_10_busy_reg;
  wire _mul_10_is_root;
  reg _mul_10_x_idle;
  reg [33-1:0] _mul_10_x_source_count;
  reg [5-1:0] _mul_10_x_source_mode;
  reg [16-1:0] _mul_10_x_source_generator_id;
  reg [32-1:0] _mul_10_x_source_offset;
  reg [33-1:0] _mul_10_x_source_size;
  reg [32-1:0] _mul_10_x_source_stride;
  reg [32-1:0] _mul_10_x_source_offset_buf;
  reg [33-1:0] _mul_10_x_source_size_buf;
  reg [32-1:0] _mul_10_x_source_stride_buf;
  reg [8-1:0] _mul_10_x_source_sel;
  reg [32-1:0] _mul_10_x_source_ram_raddr;
  reg _mul_10_x_source_ram_renable;
  wire [32-1:0] _mul_10_x_source_ram_rdata;
  reg _mul_10_x_source_fifo_deq;
  wire [32-1:0] _mul_10_x_source_fifo_rdata;
  reg [32-1:0] _mul_10_x_source_empty_data;
  reg _mul_10_y_idle;
  reg [33-1:0] _mul_10_y_source_count;
  reg [5-1:0] _mul_10_y_source_mode;
  reg [16-1:0] _mul_10_y_source_generator_id;
  reg [32-1:0] _mul_10_y_source_offset;
  reg [33-1:0] _mul_10_y_source_size;
  reg [32-1:0] _mul_10_y_source_stride;
  reg [32-1:0] _mul_10_y_source_offset_buf;
  reg [33-1:0] _mul_10_y_source_size_buf;
  reg [32-1:0] _mul_10_y_source_stride_buf;
  reg [8-1:0] _mul_10_y_source_sel;
  reg [32-1:0] _mul_10_y_source_ram_raddr;
  reg _mul_10_y_source_ram_renable;
  wire [32-1:0] _mul_10_y_source_ram_rdata;
  reg _mul_10_y_source_fifo_deq;
  wire [32-1:0] _mul_10_y_source_fifo_rdata;
  reg [32-1:0] _mul_10_y_source_empty_data;
  reg _mul_10_rshift_idle;
  reg [33-1:0] _mul_10_rshift_source_count;
  reg [5-1:0] _mul_10_rshift_source_mode;
  reg [16-1:0] _mul_10_rshift_source_generator_id;
  reg [32-1:0] _mul_10_rshift_source_offset;
  reg [33-1:0] _mul_10_rshift_source_size;
  reg [32-1:0] _mul_10_rshift_source_stride;
  reg [32-1:0] _mul_10_rshift_source_offset_buf;
  reg [33-1:0] _mul_10_rshift_source_size_buf;
  reg [32-1:0] _mul_10_rshift_source_stride_buf;
  reg [8-1:0] _mul_10_rshift_source_sel;
  reg [32-1:0] _mul_10_rshift_source_ram_raddr;
  reg _mul_10_rshift_source_ram_renable;
  wire [32-1:0] _mul_10_rshift_source_ram_rdata;
  reg _mul_10_rshift_source_fifo_deq;
  wire [32-1:0] _mul_10_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_10_rshift_source_empty_data;
  reg [33-1:0] _mul_10_z_sink_count;
  reg [5-1:0] _mul_10_z_sink_mode;
  reg [16-1:0] _mul_10_z_sink_generator_id;
  reg [32-1:0] _mul_10_z_sink_offset;
  reg [33-1:0] _mul_10_z_sink_size;
  reg [32-1:0] _mul_10_z_sink_stride;
  reg [32-1:0] _mul_10_z_sink_offset_buf;
  reg [33-1:0] _mul_10_z_sink_size_buf;
  reg [32-1:0] _mul_10_z_sink_stride_buf;
  reg [8-1:0] _mul_10_z_sink_sel;
  reg [32-1:0] _mul_10_z_sink_waddr;
  reg _mul_10_z_sink_wenable;
  reg [32-1:0] _mul_10_z_sink_wdata;
  reg _mul_10_z_sink_fifo_enq;
  reg [32-1:0] _mul_10_z_sink_fifo_wdata;
  reg [32-1:0] _mul_10_z_sink_immediate;
  reg _mul_11_stream_ivalid;
  wire _mul_11_stream_oready;
  wire _mul_11_stream_internal_oready;
  assign _mul_11_stream_internal_oready = 1;
  reg [32-1:0] _mul_11_fsm;
  localparam _mul_11_fsm_init = 0;
  wire _mul_11_run_flag;
  assign _mul_11_run_flag = 0;
  reg _mul_11_source_start;
  wire _mul_11_source_stop;
  reg _mul_11_source_busy;
  wire _mul_11_sink_start;
  wire _mul_11_sink_stop;
  wire _mul_11_sink_busy;
  wire _mul_11_busy;
  reg _mul_11_busy_reg;
  wire _mul_11_is_root;
  reg _mul_11_x_idle;
  reg [33-1:0] _mul_11_x_source_count;
  reg [5-1:0] _mul_11_x_source_mode;
  reg [16-1:0] _mul_11_x_source_generator_id;
  reg [32-1:0] _mul_11_x_source_offset;
  reg [33-1:0] _mul_11_x_source_size;
  reg [32-1:0] _mul_11_x_source_stride;
  reg [32-1:0] _mul_11_x_source_offset_buf;
  reg [33-1:0] _mul_11_x_source_size_buf;
  reg [32-1:0] _mul_11_x_source_stride_buf;
  reg [8-1:0] _mul_11_x_source_sel;
  reg [32-1:0] _mul_11_x_source_ram_raddr;
  reg _mul_11_x_source_ram_renable;
  wire [32-1:0] _mul_11_x_source_ram_rdata;
  reg _mul_11_x_source_fifo_deq;
  wire [32-1:0] _mul_11_x_source_fifo_rdata;
  reg [32-1:0] _mul_11_x_source_empty_data;
  reg _mul_11_y_idle;
  reg [33-1:0] _mul_11_y_source_count;
  reg [5-1:0] _mul_11_y_source_mode;
  reg [16-1:0] _mul_11_y_source_generator_id;
  reg [32-1:0] _mul_11_y_source_offset;
  reg [33-1:0] _mul_11_y_source_size;
  reg [32-1:0] _mul_11_y_source_stride;
  reg [32-1:0] _mul_11_y_source_offset_buf;
  reg [33-1:0] _mul_11_y_source_size_buf;
  reg [32-1:0] _mul_11_y_source_stride_buf;
  reg [8-1:0] _mul_11_y_source_sel;
  reg [32-1:0] _mul_11_y_source_ram_raddr;
  reg _mul_11_y_source_ram_renable;
  wire [32-1:0] _mul_11_y_source_ram_rdata;
  reg _mul_11_y_source_fifo_deq;
  wire [32-1:0] _mul_11_y_source_fifo_rdata;
  reg [32-1:0] _mul_11_y_source_empty_data;
  reg _mul_11_rshift_idle;
  reg [33-1:0] _mul_11_rshift_source_count;
  reg [5-1:0] _mul_11_rshift_source_mode;
  reg [16-1:0] _mul_11_rshift_source_generator_id;
  reg [32-1:0] _mul_11_rshift_source_offset;
  reg [33-1:0] _mul_11_rshift_source_size;
  reg [32-1:0] _mul_11_rshift_source_stride;
  reg [32-1:0] _mul_11_rshift_source_offset_buf;
  reg [33-1:0] _mul_11_rshift_source_size_buf;
  reg [32-1:0] _mul_11_rshift_source_stride_buf;
  reg [8-1:0] _mul_11_rshift_source_sel;
  reg [32-1:0] _mul_11_rshift_source_ram_raddr;
  reg _mul_11_rshift_source_ram_renable;
  wire [32-1:0] _mul_11_rshift_source_ram_rdata;
  reg _mul_11_rshift_source_fifo_deq;
  wire [32-1:0] _mul_11_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_11_rshift_source_empty_data;
  reg [33-1:0] _mul_11_z_sink_count;
  reg [5-1:0] _mul_11_z_sink_mode;
  reg [16-1:0] _mul_11_z_sink_generator_id;
  reg [32-1:0] _mul_11_z_sink_offset;
  reg [33-1:0] _mul_11_z_sink_size;
  reg [32-1:0] _mul_11_z_sink_stride;
  reg [32-1:0] _mul_11_z_sink_offset_buf;
  reg [33-1:0] _mul_11_z_sink_size_buf;
  reg [32-1:0] _mul_11_z_sink_stride_buf;
  reg [8-1:0] _mul_11_z_sink_sel;
  reg [32-1:0] _mul_11_z_sink_waddr;
  reg _mul_11_z_sink_wenable;
  reg [32-1:0] _mul_11_z_sink_wdata;
  reg _mul_11_z_sink_fifo_enq;
  reg [32-1:0] _mul_11_z_sink_fifo_wdata;
  reg [32-1:0] _mul_11_z_sink_immediate;
  reg _stream_conv2d_2_stream_ivalid;
  wire _stream_conv2d_2_stream_oready;
  wire _stream_conv2d_2_stream_internal_oready;
  assign _stream_conv2d_2_stream_oready = _stream_conv2d_2_stream_internal_oready;
  reg [32-1:0] _stream_conv2d_2_fsm;
  localparam _stream_conv2d_2_fsm_init = 0;
  wire _stream_conv2d_2_run_flag;
  reg _stream_conv2d_2_source_start;
  wire _stream_conv2d_2_source_stop;
  reg _stream_conv2d_2_source_busy;
  wire _stream_conv2d_2_sink_start;
  wire _stream_conv2d_2_sink_stop;
  wire _stream_conv2d_2_sink_busy;
  wire _stream_conv2d_2_busy;
  reg _stream_conv2d_2_busy_reg;
  wire _stream_conv2d_2_is_root;
  assign _stream_conv2d_2_is_root = 1;
  reg [4-1:0] _stream_conv2d_2_parameter_0_next_parameter_data;
  reg [2-1:0] _stream_conv2d_2_parameter_1_next_parameter_data;
  reg [2-1:0] _stream_conv2d_2_parameter_2_next_parameter_data;
  reg [9-1:0] _stream_conv2d_2_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_conv2d_2_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_conv2d_2_parameter_6_next_parameter_data;
  reg _stream_conv2d_2_source_7_idle;
  reg [33-1:0] _stream_conv2d_2_source_7_source_count;
  reg [5-1:0] _stream_conv2d_2_source_7_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_7_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_7_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_7_source_size;
  reg [32-1:0] _stream_conv2d_2_source_7_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_7_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_7_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_7_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_7_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_7_source_ram_raddr;
  reg _stream_conv2d_2_source_7_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_7_source_ram_rdata;
  reg _stream_conv2d_2_source_7_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_7_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_7_source_empty_data;
  reg [1-1:0] _stream_conv2d_2_parameter_8_next_parameter_data;
  reg _stream_conv2d_2_source_9_idle;
  reg [33-1:0] _stream_conv2d_2_source_9_source_count;
  reg [5-1:0] _stream_conv2d_2_source_9_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_9_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_9_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_9_source_size;
  reg [32-1:0] _stream_conv2d_2_source_9_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_9_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_9_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_9_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_9_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_9_source_ram_raddr;
  reg _stream_conv2d_2_source_9_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_9_source_ram_rdata;
  reg _stream_conv2d_2_source_9_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_9_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_9_source_empty_data;
  reg [1-1:0] _stream_conv2d_2_parameter_10_next_parameter_data;
  reg _stream_conv2d_2_source_11_idle;
  reg [33-1:0] _stream_conv2d_2_source_11_source_count;
  reg [5-1:0] _stream_conv2d_2_source_11_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_11_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_11_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_11_source_size;
  reg [32-1:0] _stream_conv2d_2_source_11_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_11_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_11_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_11_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_11_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_11_source_ram_raddr;
  reg _stream_conv2d_2_source_11_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_11_source_ram_rdata;
  reg _stream_conv2d_2_source_11_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_11_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_11_source_empty_data;
  reg [1-1:0] _stream_conv2d_2_parameter_12_next_parameter_data;
  reg _stream_conv2d_2_source_13_idle;
  reg [33-1:0] _stream_conv2d_2_source_13_source_count;
  reg [5-1:0] _stream_conv2d_2_source_13_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_13_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_13_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_13_source_size;
  reg [32-1:0] _stream_conv2d_2_source_13_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_13_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_13_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_13_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_13_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_13_source_ram_raddr;
  reg _stream_conv2d_2_source_13_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_13_source_ram_rdata;
  reg _stream_conv2d_2_source_13_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_13_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_13_source_empty_data;
  reg [1-1:0] _stream_conv2d_2_parameter_14_next_parameter_data;
  reg _stream_conv2d_2_source_15_idle;
  reg [33-1:0] _stream_conv2d_2_source_15_source_count;
  reg [5-1:0] _stream_conv2d_2_source_15_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_15_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_15_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_15_source_size;
  reg [32-1:0] _stream_conv2d_2_source_15_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_15_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_15_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_15_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_15_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_15_source_ram_raddr;
  reg _stream_conv2d_2_source_15_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_15_source_ram_rdata;
  reg _stream_conv2d_2_source_15_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_15_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_15_source_empty_data;
  reg [1-1:0] _stream_conv2d_2_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_conv2d_2_parameter_17_next_parameter_data;
  reg [1-1:0] _stream_conv2d_2_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_conv2d_2_parameter_19_next_parameter_data;
  reg _stream_conv2d_2_source_20_idle;
  reg [33-1:0] _stream_conv2d_2_source_20_source_count;
  reg [5-1:0] _stream_conv2d_2_source_20_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_20_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_20_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_20_source_size;
  reg [32-1:0] _stream_conv2d_2_source_20_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_20_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_20_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_20_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_20_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_20_source_ram_raddr;
  reg _stream_conv2d_2_source_20_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_20_source_ram_rdata;
  reg _stream_conv2d_2_source_20_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_20_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_20_source_empty_data;
  reg _stream_conv2d_2_source_21_idle;
  reg [33-1:0] _stream_conv2d_2_source_21_source_count;
  reg [5-1:0] _stream_conv2d_2_source_21_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_21_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_21_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_21_source_size;
  reg [32-1:0] _stream_conv2d_2_source_21_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_21_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_21_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_21_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_21_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_21_source_ram_raddr;
  reg _stream_conv2d_2_source_21_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_21_source_ram_rdata;
  reg _stream_conv2d_2_source_21_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_21_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_21_source_empty_data;
  reg _stream_conv2d_2_source_22_idle;
  reg [33-1:0] _stream_conv2d_2_source_22_source_count;
  reg [5-1:0] _stream_conv2d_2_source_22_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_22_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_22_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_22_source_size;
  reg [32-1:0] _stream_conv2d_2_source_22_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_22_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_22_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_22_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_22_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_22_source_ram_raddr;
  reg _stream_conv2d_2_source_22_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_22_source_ram_rdata;
  reg _stream_conv2d_2_source_22_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_22_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_22_source_empty_data;
  reg _stream_conv2d_2_source_23_idle;
  reg [33-1:0] _stream_conv2d_2_source_23_source_count;
  reg [5-1:0] _stream_conv2d_2_source_23_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_23_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_23_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_23_source_size;
  reg [32-1:0] _stream_conv2d_2_source_23_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_23_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_23_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_23_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_23_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_23_source_ram_raddr;
  reg _stream_conv2d_2_source_23_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_23_source_ram_rdata;
  reg _stream_conv2d_2_source_23_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_23_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_23_source_empty_data;
  reg _stream_conv2d_2_source_24_idle;
  reg [33-1:0] _stream_conv2d_2_source_24_source_count;
  reg [5-1:0] _stream_conv2d_2_source_24_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_24_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_24_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_24_source_size;
  reg [32-1:0] _stream_conv2d_2_source_24_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_24_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_24_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_24_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_24_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_24_source_ram_raddr;
  reg _stream_conv2d_2_source_24_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_24_source_ram_rdata;
  reg _stream_conv2d_2_source_24_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_24_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_24_source_empty_data;
  reg _stream_conv2d_2_source_25_idle;
  reg [33-1:0] _stream_conv2d_2_source_25_source_count;
  reg [5-1:0] _stream_conv2d_2_source_25_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_25_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_25_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_25_source_size;
  reg [32-1:0] _stream_conv2d_2_source_25_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_25_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_25_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_25_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_25_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_25_source_ram_raddr;
  reg _stream_conv2d_2_source_25_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_25_source_ram_rdata;
  reg _stream_conv2d_2_source_25_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_25_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_25_source_empty_data;
  reg _stream_conv2d_2_source_26_idle;
  reg [33-1:0] _stream_conv2d_2_source_26_source_count;
  reg [5-1:0] _stream_conv2d_2_source_26_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_26_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_26_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_26_source_size;
  reg [32-1:0] _stream_conv2d_2_source_26_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_26_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_26_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_26_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_26_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_26_source_ram_raddr;
  reg _stream_conv2d_2_source_26_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_26_source_ram_rdata;
  reg _stream_conv2d_2_source_26_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_26_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_26_source_empty_data;
  reg _stream_conv2d_2_source_27_idle;
  reg [33-1:0] _stream_conv2d_2_source_27_source_count;
  reg [5-1:0] _stream_conv2d_2_source_27_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_27_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_27_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_27_source_size;
  reg [32-1:0] _stream_conv2d_2_source_27_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_27_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_27_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_27_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_27_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_27_source_ram_raddr;
  reg _stream_conv2d_2_source_27_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_27_source_ram_rdata;
  reg _stream_conv2d_2_source_27_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_27_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_27_source_empty_data;
  reg _stream_conv2d_2_source_28_idle;
  reg [33-1:0] _stream_conv2d_2_source_28_source_count;
  reg [5-1:0] _stream_conv2d_2_source_28_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_28_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_28_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_28_source_size;
  reg [32-1:0] _stream_conv2d_2_source_28_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_28_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_28_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_28_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_28_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_28_source_ram_raddr;
  reg _stream_conv2d_2_source_28_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_28_source_ram_rdata;
  reg _stream_conv2d_2_source_28_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_28_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_28_source_empty_data;
  reg _stream_conv2d_2_source_29_idle;
  reg [33-1:0] _stream_conv2d_2_source_29_source_count;
  reg [5-1:0] _stream_conv2d_2_source_29_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_29_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_29_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_29_source_size;
  reg [32-1:0] _stream_conv2d_2_source_29_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_29_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_29_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_29_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_29_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_29_source_ram_raddr;
  reg _stream_conv2d_2_source_29_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_29_source_ram_rdata;
  reg _stream_conv2d_2_source_29_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_29_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_29_source_empty_data;
  reg _stream_conv2d_2_source_30_idle;
  reg [33-1:0] _stream_conv2d_2_source_30_source_count;
  reg [5-1:0] _stream_conv2d_2_source_30_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_30_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_30_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_30_source_size;
  reg [32-1:0] _stream_conv2d_2_source_30_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_30_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_30_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_30_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_30_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_30_source_ram_raddr;
  reg _stream_conv2d_2_source_30_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_30_source_ram_rdata;
  reg _stream_conv2d_2_source_30_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_30_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_30_source_empty_data;
  reg _stream_conv2d_2_source_31_idle;
  reg [33-1:0] _stream_conv2d_2_source_31_source_count;
  reg [5-1:0] _stream_conv2d_2_source_31_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_31_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_31_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_31_source_size;
  reg [32-1:0] _stream_conv2d_2_source_31_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_31_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_31_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_31_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_31_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_31_source_ram_raddr;
  reg _stream_conv2d_2_source_31_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_31_source_ram_rdata;
  reg _stream_conv2d_2_source_31_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_31_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_31_source_empty_data;
  reg _stream_conv2d_2_source_32_idle;
  reg [33-1:0] _stream_conv2d_2_source_32_source_count;
  reg [5-1:0] _stream_conv2d_2_source_32_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_32_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_32_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_32_source_size;
  reg [32-1:0] _stream_conv2d_2_source_32_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_32_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_32_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_32_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_32_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_32_source_ram_raddr;
  reg _stream_conv2d_2_source_32_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_32_source_ram_rdata;
  reg _stream_conv2d_2_source_32_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_32_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_32_source_empty_data;
  reg _stream_conv2d_2_source_33_idle;
  reg [33-1:0] _stream_conv2d_2_source_33_source_count;
  reg [5-1:0] _stream_conv2d_2_source_33_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_33_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_33_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_33_source_size;
  reg [32-1:0] _stream_conv2d_2_source_33_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_33_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_33_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_33_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_33_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_33_source_ram_raddr;
  reg _stream_conv2d_2_source_33_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_33_source_ram_rdata;
  reg _stream_conv2d_2_source_33_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_33_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_33_source_empty_data;
  reg _stream_conv2d_2_source_34_idle;
  reg [33-1:0] _stream_conv2d_2_source_34_source_count;
  reg [5-1:0] _stream_conv2d_2_source_34_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_34_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_34_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_34_source_size;
  reg [32-1:0] _stream_conv2d_2_source_34_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_34_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_34_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_34_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_34_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_34_source_ram_raddr;
  reg _stream_conv2d_2_source_34_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_34_source_ram_rdata;
  reg _stream_conv2d_2_source_34_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_34_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_34_source_empty_data;
  reg _stream_conv2d_2_source_35_idle;
  reg [33-1:0] _stream_conv2d_2_source_35_source_count;
  reg [5-1:0] _stream_conv2d_2_source_35_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_35_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_35_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_35_source_size;
  reg [32-1:0] _stream_conv2d_2_source_35_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_35_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_35_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_35_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_35_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_35_source_ram_raddr;
  reg _stream_conv2d_2_source_35_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_35_source_ram_rdata;
  reg _stream_conv2d_2_source_35_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_35_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_35_source_empty_data;
  reg _stream_conv2d_2_source_36_idle;
  reg [33-1:0] _stream_conv2d_2_source_36_source_count;
  reg [5-1:0] _stream_conv2d_2_source_36_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_36_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_36_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_36_source_size;
  reg [32-1:0] _stream_conv2d_2_source_36_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_36_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_36_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_36_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_36_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_36_source_ram_raddr;
  reg _stream_conv2d_2_source_36_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_36_source_ram_rdata;
  reg _stream_conv2d_2_source_36_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_36_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_36_source_empty_data;
  reg _stream_conv2d_2_source_37_idle;
  reg [33-1:0] _stream_conv2d_2_source_37_source_count;
  reg [5-1:0] _stream_conv2d_2_source_37_source_mode;
  reg [16-1:0] _stream_conv2d_2_source_37_source_generator_id;
  reg [32-1:0] _stream_conv2d_2_source_37_source_offset;
  reg [33-1:0] _stream_conv2d_2_source_37_source_size;
  reg [32-1:0] _stream_conv2d_2_source_37_source_stride;
  reg [32-1:0] _stream_conv2d_2_source_37_source_offset_buf;
  reg [33-1:0] _stream_conv2d_2_source_37_source_size_buf;
  reg [32-1:0] _stream_conv2d_2_source_37_source_stride_buf;
  reg [8-1:0] _stream_conv2d_2_source_37_source_sel;
  reg [32-1:0] _stream_conv2d_2_source_37_source_ram_raddr;
  reg _stream_conv2d_2_source_37_source_ram_renable;
  wire [32-1:0] _stream_conv2d_2_source_37_source_ram_rdata;
  reg _stream_conv2d_2_source_37_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_2_source_37_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_2_source_37_source_empty_data;
  wire signed [32-1:0] mul_3_x_data;
  wire signed [32-1:0] mul_3_y_data;
  wire [6-1:0] mul_3_rshift_data;
  reg __mul_3_stream_ivalid_1;
  reg __mul_3_stream_ivalid_2;
  reg __mul_3_stream_ivalid_3;
  reg __mul_3_stream_ivalid_4;
  reg __mul_3_stream_ivalid_5;
  reg __mul_3_stream_ivalid_6;
  reg __mul_3_stream_ivalid_7;
  reg __mul_3_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_73;
  reg [6-1:0] _minus_data_75;
  reg [1-1:0] _greatereq_data_86;
  reg signed [32-1:0] __delay_data_641__variable_70;
  reg signed [32-1:0] __delay_data_644__variable_71;
  reg [6-1:0] __delay_data_647__variable_72;
  reg signed [66-1:0] _sll_data_77;
  reg [1-1:0] __delay_data_638_greaterthan_73;
  reg [1-1:0] __delay_data_639_greatereq_86;
  reg signed [32-1:0] __delay_data_642__delay_641__variable_70;
  reg signed [32-1:0] __delay_data_645__delay_644__variable_71;
  reg [6-1:0] __delay_data_648__delay_647__variable_72;
  reg signed [32-1:0] _cond_data_83;
  reg [1-1:0] __delay_data_640__delay_639_greatereq_86;
  reg signed [32-1:0] __delay_data_643__delay_642__delay_641__variable_70;
  reg signed [32-1:0] __delay_data_646__delay_645__delay_644__variable_71;
  reg [6-1:0] __delay_data_649__delay_648__delay_647__variable_72;
  wire signed [32-1:0] _uminus_data_85;
  assign _uminus_data_85 = -_cond_data_83;
  wire signed [32-1:0] _cond_data_88;
  assign _cond_data_88 = (__delay_data_640__delay_639_greatereq_86)? _cond_data_83 : _uminus_data_85;
  wire signed [64-1:0] __muladd_madd_odata_89;
  reg signed [64-1:0] __muladd_madd_odata_reg_89;
  wire signed [32-1:0] __muladd_data_89;
  assign __muladd_data_89 = __muladd_madd_odata_reg_89;
  wire __muladd_madd_update_89;
  assign __muladd_madd_update_89 = _mul_3_stream_oready;

  madd_0
  __muladd_madd_89
  (
    .CLK(CLK),
    .update(__muladd_madd_update_89),
    .a(__delay_data_643__delay_642__delay_641__variable_70),
    .b(__delay_data_646__delay_645__delay_644__variable_71),
    .c(_cond_data_88),
    .d(__muladd_madd_odata_89)
  );

  reg [6-1:0] __delay_data_650__delay_649__delay_648__delay_647__variable_72;
  reg [6-1:0] __delay_data_651__delay_650__delay_649__delay_648____variable_72;
  reg [6-1:0] __delay_data_652__delay_651__delay_650__delay_649____variable_72;
  reg [6-1:0] __delay_data_653__delay_652__delay_651__delay_650____variable_72;
  reg signed [32-1:0] _sra_data_90;
  wire signed [32-1:0] mul_3_z_data;
  assign mul_3_z_data = _sra_data_90;
  wire signed [32-1:0] mul_4_x_data;
  wire signed [32-1:0] mul_4_y_data;
  wire [6-1:0] mul_4_rshift_data;
  reg __mul_4_stream_ivalid_1;
  reg __mul_4_stream_ivalid_2;
  reg __mul_4_stream_ivalid_3;
  reg __mul_4_stream_ivalid_4;
  reg __mul_4_stream_ivalid_5;
  reg __mul_4_stream_ivalid_6;
  reg __mul_4_stream_ivalid_7;
  reg __mul_4_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_94;
  reg [6-1:0] _minus_data_96;
  reg [1-1:0] _greatereq_data_107;
  reg signed [32-1:0] __delay_data_660__variable_91;
  reg signed [32-1:0] __delay_data_663__variable_92;
  reg [6-1:0] __delay_data_666__variable_93;
  reg signed [66-1:0] _sll_data_98;
  reg [1-1:0] __delay_data_657_greaterthan_94;
  reg [1-1:0] __delay_data_658_greatereq_107;
  reg signed [32-1:0] __delay_data_661__delay_660__variable_91;
  reg signed [32-1:0] __delay_data_664__delay_663__variable_92;
  reg [6-1:0] __delay_data_667__delay_666__variable_93;
  reg signed [32-1:0] _cond_data_104;
  reg [1-1:0] __delay_data_659__delay_658_greatereq_107;
  reg signed [32-1:0] __delay_data_662__delay_661__delay_660__variable_91;
  reg signed [32-1:0] __delay_data_665__delay_664__delay_663__variable_92;
  reg [6-1:0] __delay_data_668__delay_667__delay_666__variable_93;
  wire signed [32-1:0] _uminus_data_106;
  assign _uminus_data_106 = -_cond_data_104;
  wire signed [32-1:0] _cond_data_109;
  assign _cond_data_109 = (__delay_data_659__delay_658_greatereq_107)? _cond_data_104 : _uminus_data_106;
  wire signed [64-1:0] __muladd_madd_odata_110;
  reg signed [64-1:0] __muladd_madd_odata_reg_110;
  wire signed [32-1:0] __muladd_data_110;
  assign __muladd_data_110 = __muladd_madd_odata_reg_110;
  wire __muladd_madd_update_110;
  assign __muladd_madd_update_110 = _mul_4_stream_oready;

  madd_1
  __muladd_madd_110
  (
    .CLK(CLK),
    .update(__muladd_madd_update_110),
    .a(__delay_data_662__delay_661__delay_660__variable_91),
    .b(__delay_data_665__delay_664__delay_663__variable_92),
    .c(_cond_data_109),
    .d(__muladd_madd_odata_110)
  );

  reg [6-1:0] __delay_data_669__delay_668__delay_667__delay_666__variable_93;
  reg [6-1:0] __delay_data_670__delay_669__delay_668__delay_667____variable_93;
  reg [6-1:0] __delay_data_671__delay_670__delay_669__delay_668____variable_93;
  reg [6-1:0] __delay_data_672__delay_671__delay_670__delay_669____variable_93;
  reg signed [32-1:0] _sra_data_111;
  wire signed [32-1:0] mul_4_z_data;
  assign mul_4_z_data = _sra_data_111;
  wire signed [32-1:0] mul_5_x_data;
  wire signed [32-1:0] mul_5_y_data;
  wire [6-1:0] mul_5_rshift_data;
  reg __mul_5_stream_ivalid_1;
  reg __mul_5_stream_ivalid_2;
  reg __mul_5_stream_ivalid_3;
  reg __mul_5_stream_ivalid_4;
  reg __mul_5_stream_ivalid_5;
  reg __mul_5_stream_ivalid_6;
  reg __mul_5_stream_ivalid_7;
  reg __mul_5_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_115;
  reg [6-1:0] _minus_data_117;
  reg [1-1:0] _greatereq_data_128;
  reg signed [32-1:0] __delay_data_679__variable_112;
  reg signed [32-1:0] __delay_data_682__variable_113;
  reg [6-1:0] __delay_data_685__variable_114;
  reg signed [66-1:0] _sll_data_119;
  reg [1-1:0] __delay_data_676_greaterthan_115;
  reg [1-1:0] __delay_data_677_greatereq_128;
  reg signed [32-1:0] __delay_data_680__delay_679__variable_112;
  reg signed [32-1:0] __delay_data_683__delay_682__variable_113;
  reg [6-1:0] __delay_data_686__delay_685__variable_114;
  reg signed [32-1:0] _cond_data_125;
  reg [1-1:0] __delay_data_678__delay_677_greatereq_128;
  reg signed [32-1:0] __delay_data_681__delay_680__delay_679__variable_112;
  reg signed [32-1:0] __delay_data_684__delay_683__delay_682__variable_113;
  reg [6-1:0] __delay_data_687__delay_686__delay_685__variable_114;
  wire signed [32-1:0] _uminus_data_127;
  assign _uminus_data_127 = -_cond_data_125;
  wire signed [32-1:0] _cond_data_130;
  assign _cond_data_130 = (__delay_data_678__delay_677_greatereq_128)? _cond_data_125 : _uminus_data_127;
  wire signed [64-1:0] __muladd_madd_odata_131;
  reg signed [64-1:0] __muladd_madd_odata_reg_131;
  wire signed [32-1:0] __muladd_data_131;
  assign __muladd_data_131 = __muladd_madd_odata_reg_131;
  wire __muladd_madd_update_131;
  assign __muladd_madd_update_131 = _mul_5_stream_oready;

  madd_2
  __muladd_madd_131
  (
    .CLK(CLK),
    .update(__muladd_madd_update_131),
    .a(__delay_data_681__delay_680__delay_679__variable_112),
    .b(__delay_data_684__delay_683__delay_682__variable_113),
    .c(_cond_data_130),
    .d(__muladd_madd_odata_131)
  );

  reg [6-1:0] __delay_data_688__delay_687__delay_686____variable_114;
  reg [6-1:0] __delay_data_689__delay_688__delay_687____variable_114;
  reg [6-1:0] __delay_data_690__delay_689__delay_688____variable_114;
  reg [6-1:0] __delay_data_691__delay_690__delay_689____variable_114;
  reg signed [32-1:0] _sra_data_132;
  wire signed [32-1:0] mul_5_z_data;
  assign mul_5_z_data = _sra_data_132;
  wire signed [32-1:0] mul_6_x_data;
  wire signed [32-1:0] mul_6_y_data;
  wire [6-1:0] mul_6_rshift_data;
  reg __mul_6_stream_ivalid_1;
  reg __mul_6_stream_ivalid_2;
  reg __mul_6_stream_ivalid_3;
  reg __mul_6_stream_ivalid_4;
  reg __mul_6_stream_ivalid_5;
  reg __mul_6_stream_ivalid_6;
  reg __mul_6_stream_ivalid_7;
  reg __mul_6_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_136;
  reg [6-1:0] _minus_data_138;
  reg [1-1:0] _greatereq_data_149;
  reg signed [32-1:0] __delay_data_698__variable_133;
  reg signed [32-1:0] __delay_data_701__variable_134;
  reg [6-1:0] __delay_data_704__variable_135;
  reg signed [66-1:0] _sll_data_140;
  reg [1-1:0] __delay_data_695_greaterthan_136;
  reg [1-1:0] __delay_data_696_greatereq_149;
  reg signed [32-1:0] __delay_data_699__delay_698__variable_133;
  reg signed [32-1:0] __delay_data_702__delay_701__variable_134;
  reg [6-1:0] __delay_data_705__delay_704__variable_135;
  reg signed [32-1:0] _cond_data_146;
  reg [1-1:0] __delay_data_697__delay_696_greatereq_149;
  reg signed [32-1:0] __delay_data_700__delay_699__delay_698__variable_133;
  reg signed [32-1:0] __delay_data_703__delay_702__delay_701__variable_134;
  reg [6-1:0] __delay_data_706__delay_705__delay_704__variable_135;
  wire signed [32-1:0] _uminus_data_148;
  assign _uminus_data_148 = -_cond_data_146;
  wire signed [32-1:0] _cond_data_151;
  assign _cond_data_151 = (__delay_data_697__delay_696_greatereq_149)? _cond_data_146 : _uminus_data_148;
  wire signed [64-1:0] __muladd_madd_odata_152;
  reg signed [64-1:0] __muladd_madd_odata_reg_152;
  wire signed [32-1:0] __muladd_data_152;
  assign __muladd_data_152 = __muladd_madd_odata_reg_152;
  wire __muladd_madd_update_152;
  assign __muladd_madd_update_152 = _mul_6_stream_oready;

  madd_3
  __muladd_madd_152
  (
    .CLK(CLK),
    .update(__muladd_madd_update_152),
    .a(__delay_data_700__delay_699__delay_698__variable_133),
    .b(__delay_data_703__delay_702__delay_701__variable_134),
    .c(_cond_data_151),
    .d(__muladd_madd_odata_152)
  );

  reg [6-1:0] __delay_data_707__delay_706__delay_705____variable_135;
  reg [6-1:0] __delay_data_708__delay_707__delay_706____variable_135;
  reg [6-1:0] __delay_data_709__delay_708__delay_707____variable_135;
  reg [6-1:0] __delay_data_710__delay_709__delay_708____variable_135;
  reg signed [32-1:0] _sra_data_153;
  wire signed [32-1:0] mul_6_z_data;
  assign mul_6_z_data = _sra_data_153;
  wire signed [32-1:0] mul_7_x_data;
  wire signed [32-1:0] mul_7_y_data;
  wire [6-1:0] mul_7_rshift_data;
  reg __mul_7_stream_ivalid_1;
  reg __mul_7_stream_ivalid_2;
  reg __mul_7_stream_ivalid_3;
  reg __mul_7_stream_ivalid_4;
  reg __mul_7_stream_ivalid_5;
  reg __mul_7_stream_ivalid_6;
  reg __mul_7_stream_ivalid_7;
  reg __mul_7_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_157;
  reg [6-1:0] _minus_data_159;
  reg [1-1:0] _greatereq_data_170;
  reg signed [32-1:0] __delay_data_717__variable_154;
  reg signed [32-1:0] __delay_data_720__variable_155;
  reg [6-1:0] __delay_data_723__variable_156;
  reg signed [66-1:0] _sll_data_161;
  reg [1-1:0] __delay_data_714_greaterthan_157;
  reg [1-1:0] __delay_data_715_greatereq_170;
  reg signed [32-1:0] __delay_data_718__delay_717__variable_154;
  reg signed [32-1:0] __delay_data_721__delay_720__variable_155;
  reg [6-1:0] __delay_data_724__delay_723__variable_156;
  reg signed [32-1:0] _cond_data_167;
  reg [1-1:0] __delay_data_716__delay_715_greatereq_170;
  reg signed [32-1:0] __delay_data_719__delay_718__delay_717__variable_154;
  reg signed [32-1:0] __delay_data_722__delay_721__delay_720__variable_155;
  reg [6-1:0] __delay_data_725__delay_724__delay_723__variable_156;
  wire signed [32-1:0] _uminus_data_169;
  assign _uminus_data_169 = -_cond_data_167;
  wire signed [32-1:0] _cond_data_172;
  assign _cond_data_172 = (__delay_data_716__delay_715_greatereq_170)? _cond_data_167 : _uminus_data_169;
  wire signed [64-1:0] __muladd_madd_odata_173;
  reg signed [64-1:0] __muladd_madd_odata_reg_173;
  wire signed [32-1:0] __muladd_data_173;
  assign __muladd_data_173 = __muladd_madd_odata_reg_173;
  wire __muladd_madd_update_173;
  assign __muladd_madd_update_173 = _mul_7_stream_oready;

  madd_4
  __muladd_madd_173
  (
    .CLK(CLK),
    .update(__muladd_madd_update_173),
    .a(__delay_data_719__delay_718__delay_717__variable_154),
    .b(__delay_data_722__delay_721__delay_720__variable_155),
    .c(_cond_data_172),
    .d(__muladd_madd_odata_173)
  );

  reg [6-1:0] __delay_data_726__delay_725__delay_724____variable_156;
  reg [6-1:0] __delay_data_727__delay_726__delay_725____variable_156;
  reg [6-1:0] __delay_data_728__delay_727__delay_726____variable_156;
  reg [6-1:0] __delay_data_729__delay_728__delay_727____variable_156;
  reg signed [32-1:0] _sra_data_174;
  wire signed [32-1:0] mul_7_z_data;
  assign mul_7_z_data = _sra_data_174;
  wire signed [32-1:0] mul_8_x_data;
  wire signed [32-1:0] mul_8_y_data;
  wire [6-1:0] mul_8_rshift_data;
  reg __mul_8_stream_ivalid_1;
  reg __mul_8_stream_ivalid_2;
  reg __mul_8_stream_ivalid_3;
  reg __mul_8_stream_ivalid_4;
  reg __mul_8_stream_ivalid_5;
  reg __mul_8_stream_ivalid_6;
  reg __mul_8_stream_ivalid_7;
  reg __mul_8_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_178;
  reg [6-1:0] _minus_data_180;
  reg [1-1:0] _greatereq_data_191;
  reg signed [32-1:0] __delay_data_736__variable_175;
  reg signed [32-1:0] __delay_data_739__variable_176;
  reg [6-1:0] __delay_data_742__variable_177;
  reg signed [66-1:0] _sll_data_182;
  reg [1-1:0] __delay_data_733_greaterthan_178;
  reg [1-1:0] __delay_data_734_greatereq_191;
  reg signed [32-1:0] __delay_data_737__delay_736__variable_175;
  reg signed [32-1:0] __delay_data_740__delay_739__variable_176;
  reg [6-1:0] __delay_data_743__delay_742__variable_177;
  reg signed [32-1:0] _cond_data_188;
  reg [1-1:0] __delay_data_735__delay_734_greatereq_191;
  reg signed [32-1:0] __delay_data_738__delay_737__delay_736__variable_175;
  reg signed [32-1:0] __delay_data_741__delay_740__delay_739__variable_176;
  reg [6-1:0] __delay_data_744__delay_743__delay_742__variable_177;
  wire signed [32-1:0] _uminus_data_190;
  assign _uminus_data_190 = -_cond_data_188;
  wire signed [32-1:0] _cond_data_193;
  assign _cond_data_193 = (__delay_data_735__delay_734_greatereq_191)? _cond_data_188 : _uminus_data_190;
  wire signed [64-1:0] __muladd_madd_odata_194;
  reg signed [64-1:0] __muladd_madd_odata_reg_194;
  wire signed [32-1:0] __muladd_data_194;
  assign __muladd_data_194 = __muladd_madd_odata_reg_194;
  wire __muladd_madd_update_194;
  assign __muladd_madd_update_194 = _mul_8_stream_oready;

  madd_5
  __muladd_madd_194
  (
    .CLK(CLK),
    .update(__muladd_madd_update_194),
    .a(__delay_data_738__delay_737__delay_736__variable_175),
    .b(__delay_data_741__delay_740__delay_739__variable_176),
    .c(_cond_data_193),
    .d(__muladd_madd_odata_194)
  );

  reg [6-1:0] __delay_data_745__delay_744__delay_743____variable_177;
  reg [6-1:0] __delay_data_746__delay_745__delay_744____variable_177;
  reg [6-1:0] __delay_data_747__delay_746__delay_745____variable_177;
  reg [6-1:0] __delay_data_748__delay_747__delay_746____variable_177;
  reg signed [32-1:0] _sra_data_195;
  wire signed [32-1:0] mul_8_z_data;
  assign mul_8_z_data = _sra_data_195;
  wire signed [32-1:0] mul_9_x_data;
  wire signed [32-1:0] mul_9_y_data;
  wire [6-1:0] mul_9_rshift_data;
  reg __mul_9_stream_ivalid_1;
  reg __mul_9_stream_ivalid_2;
  reg __mul_9_stream_ivalid_3;
  reg __mul_9_stream_ivalid_4;
  reg __mul_9_stream_ivalid_5;
  reg __mul_9_stream_ivalid_6;
  reg __mul_9_stream_ivalid_7;
  reg __mul_9_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_199;
  reg [6-1:0] _minus_data_201;
  reg [1-1:0] _greatereq_data_212;
  reg signed [32-1:0] __delay_data_755__variable_196;
  reg signed [32-1:0] __delay_data_758__variable_197;
  reg [6-1:0] __delay_data_761__variable_198;
  reg signed [66-1:0] _sll_data_203;
  reg [1-1:0] __delay_data_752_greaterthan_199;
  reg [1-1:0] __delay_data_753_greatereq_212;
  reg signed [32-1:0] __delay_data_756__delay_755__variable_196;
  reg signed [32-1:0] __delay_data_759__delay_758__variable_197;
  reg [6-1:0] __delay_data_762__delay_761__variable_198;
  reg signed [32-1:0] _cond_data_209;
  reg [1-1:0] __delay_data_754__delay_753_greatereq_212;
  reg signed [32-1:0] __delay_data_757__delay_756__delay_755__variable_196;
  reg signed [32-1:0] __delay_data_760__delay_759__delay_758__variable_197;
  reg [6-1:0] __delay_data_763__delay_762__delay_761__variable_198;
  wire signed [32-1:0] _uminus_data_211;
  assign _uminus_data_211 = -_cond_data_209;
  wire signed [32-1:0] _cond_data_214;
  assign _cond_data_214 = (__delay_data_754__delay_753_greatereq_212)? _cond_data_209 : _uminus_data_211;
  wire signed [64-1:0] __muladd_madd_odata_215;
  reg signed [64-1:0] __muladd_madd_odata_reg_215;
  wire signed [32-1:0] __muladd_data_215;
  assign __muladd_data_215 = __muladd_madd_odata_reg_215;
  wire __muladd_madd_update_215;
  assign __muladd_madd_update_215 = _mul_9_stream_oready;

  madd_6
  __muladd_madd_215
  (
    .CLK(CLK),
    .update(__muladd_madd_update_215),
    .a(__delay_data_757__delay_756__delay_755__variable_196),
    .b(__delay_data_760__delay_759__delay_758__variable_197),
    .c(_cond_data_214),
    .d(__muladd_madd_odata_215)
  );

  reg [6-1:0] __delay_data_764__delay_763__delay_762____variable_198;
  reg [6-1:0] __delay_data_765__delay_764__delay_763____variable_198;
  reg [6-1:0] __delay_data_766__delay_765__delay_764____variable_198;
  reg [6-1:0] __delay_data_767__delay_766__delay_765____variable_198;
  reg signed [32-1:0] _sra_data_216;
  wire signed [32-1:0] mul_9_z_data;
  assign mul_9_z_data = _sra_data_216;
  wire signed [32-1:0] mul_10_x_data;
  wire signed [32-1:0] mul_10_y_data;
  wire [6-1:0] mul_10_rshift_data;
  reg __mul_10_stream_ivalid_1;
  reg __mul_10_stream_ivalid_2;
  reg __mul_10_stream_ivalid_3;
  reg __mul_10_stream_ivalid_4;
  reg __mul_10_stream_ivalid_5;
  reg __mul_10_stream_ivalid_6;
  reg __mul_10_stream_ivalid_7;
  reg __mul_10_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_220;
  reg [6-1:0] _minus_data_222;
  reg [1-1:0] _greatereq_data_233;
  reg signed [32-1:0] __delay_data_774__variable_217;
  reg signed [32-1:0] __delay_data_777__variable_218;
  reg [6-1:0] __delay_data_780__variable_219;
  reg signed [66-1:0] _sll_data_224;
  reg [1-1:0] __delay_data_771_greaterthan_220;
  reg [1-1:0] __delay_data_772_greatereq_233;
  reg signed [32-1:0] __delay_data_775__delay_774__variable_217;
  reg signed [32-1:0] __delay_data_778__delay_777__variable_218;
  reg [6-1:0] __delay_data_781__delay_780__variable_219;
  reg signed [32-1:0] _cond_data_230;
  reg [1-1:0] __delay_data_773__delay_772_greatereq_233;
  reg signed [32-1:0] __delay_data_776__delay_775__delay_774__variable_217;
  reg signed [32-1:0] __delay_data_779__delay_778__delay_777__variable_218;
  reg [6-1:0] __delay_data_782__delay_781__delay_780__variable_219;
  wire signed [32-1:0] _uminus_data_232;
  assign _uminus_data_232 = -_cond_data_230;
  wire signed [32-1:0] _cond_data_235;
  assign _cond_data_235 = (__delay_data_773__delay_772_greatereq_233)? _cond_data_230 : _uminus_data_232;
  wire signed [64-1:0] __muladd_madd_odata_236;
  reg signed [64-1:0] __muladd_madd_odata_reg_236;
  wire signed [32-1:0] __muladd_data_236;
  assign __muladd_data_236 = __muladd_madd_odata_reg_236;
  wire __muladd_madd_update_236;
  assign __muladd_madd_update_236 = _mul_10_stream_oready;

  madd_7
  __muladd_madd_236
  (
    .CLK(CLK),
    .update(__muladd_madd_update_236),
    .a(__delay_data_776__delay_775__delay_774__variable_217),
    .b(__delay_data_779__delay_778__delay_777__variable_218),
    .c(_cond_data_235),
    .d(__muladd_madd_odata_236)
  );

  reg [6-1:0] __delay_data_783__delay_782__delay_781____variable_219;
  reg [6-1:0] __delay_data_784__delay_783__delay_782____variable_219;
  reg [6-1:0] __delay_data_785__delay_784__delay_783____variable_219;
  reg [6-1:0] __delay_data_786__delay_785__delay_784____variable_219;
  reg signed [32-1:0] _sra_data_237;
  wire signed [32-1:0] mul_10_z_data;
  assign mul_10_z_data = _sra_data_237;
  wire signed [32-1:0] mul_11_x_data;
  wire signed [32-1:0] mul_11_y_data;
  wire [6-1:0] mul_11_rshift_data;
  reg __mul_11_stream_ivalid_1;
  reg __mul_11_stream_ivalid_2;
  reg __mul_11_stream_ivalid_3;
  reg __mul_11_stream_ivalid_4;
  reg __mul_11_stream_ivalid_5;
  reg __mul_11_stream_ivalid_6;
  reg __mul_11_stream_ivalid_7;
  reg __mul_11_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_241;
  reg [6-1:0] _minus_data_243;
  reg [1-1:0] _greatereq_data_254;
  reg signed [32-1:0] __delay_data_793__variable_238;
  reg signed [32-1:0] __delay_data_796__variable_239;
  reg [6-1:0] __delay_data_799__variable_240;
  reg signed [66-1:0] _sll_data_245;
  reg [1-1:0] __delay_data_790_greaterthan_241;
  reg [1-1:0] __delay_data_791_greatereq_254;
  reg signed [32-1:0] __delay_data_794__delay_793__variable_238;
  reg signed [32-1:0] __delay_data_797__delay_796__variable_239;
  reg [6-1:0] __delay_data_800__delay_799__variable_240;
  reg signed [32-1:0] _cond_data_251;
  reg [1-1:0] __delay_data_792__delay_791_greatereq_254;
  reg signed [32-1:0] __delay_data_795__delay_794__delay_793__variable_238;
  reg signed [32-1:0] __delay_data_798__delay_797__delay_796__variable_239;
  reg [6-1:0] __delay_data_801__delay_800__delay_799__variable_240;
  wire signed [32-1:0] _uminus_data_253;
  assign _uminus_data_253 = -_cond_data_251;
  wire signed [32-1:0] _cond_data_256;
  assign _cond_data_256 = (__delay_data_792__delay_791_greatereq_254)? _cond_data_251 : _uminus_data_253;
  wire signed [64-1:0] __muladd_madd_odata_257;
  reg signed [64-1:0] __muladd_madd_odata_reg_257;
  wire signed [32-1:0] __muladd_data_257;
  assign __muladd_data_257 = __muladd_madd_odata_reg_257;
  wire __muladd_madd_update_257;
  assign __muladd_madd_update_257 = _mul_11_stream_oready;

  madd_8
  __muladd_madd_257
  (
    .CLK(CLK),
    .update(__muladd_madd_update_257),
    .a(__delay_data_795__delay_794__delay_793__variable_238),
    .b(__delay_data_798__delay_797__delay_796__variable_239),
    .c(_cond_data_256),
    .d(__muladd_madd_odata_257)
  );

  reg [6-1:0] __delay_data_802__delay_801__delay_800____variable_240;
  reg [6-1:0] __delay_data_803__delay_802__delay_801____variable_240;
  reg [6-1:0] __delay_data_804__delay_803__delay_802____variable_240;
  reg [6-1:0] __delay_data_805__delay_804__delay_803____variable_240;
  reg signed [32-1:0] _sra_data_258;
  wire signed [32-1:0] mul_11_z_data;
  assign mul_11_z_data = _sra_data_258;
  wire signed [32-1:0] add_tree_1_var0_data;
  wire signed [32-1:0] add_tree_1_var1_data;
  wire signed [32-1:0] add_tree_1_var2_data;
  wire signed [32-1:0] add_tree_1_var3_data;
  wire signed [32-1:0] add_tree_1_var4_data;
  wire signed [32-1:0] add_tree_1_var5_data;
  wire signed [32-1:0] add_tree_1_var6_data;
  wire signed [32-1:0] add_tree_1_var7_data;
  wire signed [32-1:0] add_tree_1_var8_data;
  reg __add_tree_1_stream_ivalid_1;
  reg __add_tree_1_stream_ivalid_2;
  reg signed [32-1:0] __plusn_data_32;
  reg signed [32-1:0] __plusn_data_33;
  reg signed [32-1:0] __plusn_data_34;
  reg signed [32-1:0] __plusn_data_35;
  wire signed [32-1:0] add_tree_1_sum_data;
  assign add_tree_1_sum_data = __plusn_data_35;
  wire signed [32-1:0] acc_0_x_data;
  wire [6-1:0] acc_0_rshift_data;
  wire [32-1:0] acc_0_size_data;
  wire [1-1:0] acc_0__reduce_reset_data;
  reg __acc_0_stream_ivalid_1;
  reg __acc_0_stream_ivalid_2;
  reg __acc_0_stream_ivalid_3;
  reg __acc_0_stream_ivalid_4;
  reg __acc_0_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_3;
  reg [6-1:0] _minus_data_5;
  reg signed [32-1:0] _reduceadd_data_16;
  reg [33-1:0] _reduceadd_count_16;
  reg _reduceadd_prev_count_max_16;
  wire _reduceadd_reset_cond_16;
  assign _reduceadd_reset_cond_16 = acc_0__reduce_reset_data || _reduceadd_prev_count_max_16;
  wire [33-1:0] _reduceadd_current_count_16;
  assign _reduceadd_current_count_16 = (_reduceadd_reset_cond_16)? 0 : _reduceadd_count_16;
  wire signed [32-1:0] _reduceadd_current_data_16;
  assign _reduceadd_current_data_16 = (_reduceadd_reset_cond_16)? 1'sd0 : _reduceadd_data_16;
  reg [1-1:0] _pulse_data_18;
  reg [33-1:0] _pulse_count_18;
  reg _pulse_prev_count_max_18;
  wire _pulse_reset_cond_18;
  assign _pulse_reset_cond_18 = acc_0__reduce_reset_data || _pulse_prev_count_max_18;
  wire [33-1:0] _pulse_current_count_18;
  assign _pulse_current_count_18 = (_pulse_reset_cond_18)? 0 : _pulse_count_18;
  wire [1-1:0] _pulse_current_data_18;
  assign _pulse_current_data_18 = (_pulse_reset_cond_18)? 1'sd0 : _pulse_data_18;
  reg [6-1:0] __delay_data_814__variable_1;
  reg signed [66-1:0] _sll_data_7;
  reg [1-1:0] __delay_data_811_greaterthan_3;
  reg signed [32-1:0] __delay_data_812_reduceadd_16;
  reg [6-1:0] __delay_data_815__delay_814__variable_1;
  reg [1-1:0] __delay_data_818_pulse_18;
  reg signed [32-1:0] _cond_data_13;
  reg signed [32-1:0] __delay_data_813__delay_812_reduceadd_16;
  reg [6-1:0] __delay_data_816__delay_815__delay_814__variable_1;
  reg [1-1:0] __delay_data_819__delay_818_pulse_18;
  reg signed [32-1:0] _plus_data_20;
  reg [6-1:0] __delay_data_817__delay_816__delay_815__delay_814__variable_1;
  reg [1-1:0] __delay_data_820__delay_819__delay_818_pulse_18;
  reg signed [32-1:0] _sra_data_21;
  reg [1-1:0] __delay_data_821__delay_820__delay_819__delay_818_pulse_18;
  wire signed [32-1:0] acc_0_sum_data;
  assign acc_0_sum_data = _sra_data_21;
  wire [1-1:0] acc_0_valid_data;
  assign acc_0_valid_data = __delay_data_821__delay_820__delay_819__delay_818_pulse_18;
  wire signed [32-1:0] mul_rshift_round_clip_2_x_data;
  wire signed [32-1:0] mul_rshift_round_clip_2_y_data;
  wire [6-1:0] mul_rshift_round_clip_2_rshift_data;
  reg __mul_rshift_round_clip_2_stream_ivalid_1;
  reg __mul_rshift_round_clip_2_stream_ivalid_2;
  reg __mul_rshift_round_clip_2_stream_ivalid_3;
  reg __mul_rshift_round_clip_2_stream_ivalid_4;
  reg __mul_rshift_round_clip_2_stream_ivalid_5;
  reg __mul_rshift_round_clip_2_stream_ivalid_6;
  reg __mul_rshift_round_clip_2_stream_ivalid_7;
  reg __mul_rshift_round_clip_2_stream_ivalid_8;
  wire signed [64-1:0] _times_mul_odata_39;
  reg signed [64-1:0] _times_mul_odata_reg_39;
  wire signed [64-1:0] _times_data_39;
  assign _times_data_39 = _times_mul_odata_reg_39;
  wire _times_mul_update_39;
  assign _times_mul_update_39 = _mul_rshift_round_clip_2_stream_oready;

  multiplier_0
  _times_mul_39
  (
    .CLK(CLK),
    .update(_times_mul_update_39),
    .a(mul_rshift_round_clip_2_x_data),
    .b(mul_rshift_round_clip_2_y_data),
    .c(_times_mul_odata_39)
  );

  wire [6-1:0] _minus_data_42;
  assign _minus_data_42 = mul_rshift_round_clip_2_rshift_data - 2'sd1;
  wire signed [66-1:0] _sll_data_45;
  assign _sll_data_45 = 2'sd1 << _minus_data_42;
  wire [1-1:0] _eq_data_57;
  assign _eq_data_57 = mul_rshift_round_clip_2_rshift_data == 1'sd0;
  reg signed [66-1:0] __delay_data_827_sll_45;
  reg [6-1:0] __delay_data_831__variable_38;
  reg [1-1:0] __delay_data_835_eq_57;
  reg signed [66-1:0] __delay_data_828__delay_827_sll_45;
  reg [6-1:0] __delay_data_832__delay_831__variable_38;
  reg [1-1:0] __delay_data_836__delay_835_eq_57;
  reg signed [66-1:0] __delay_data_829__delay_828__delay_827_sll_45;
  reg [6-1:0] __delay_data_833__delay_832__delay_831__variable_38;
  reg [1-1:0] __delay_data_837__delay_836__delay_835_eq_57;
  reg signed [66-1:0] __delay_data_830__delay_829__delay_828__delay_827_sll_45;
  reg [6-1:0] __delay_data_834__delay_833__delay_832__delay_831__variable_38;
  reg [1-1:0] __delay_data_838__delay_837__delay_836__delay_835_eq_57;
  wire [1-1:0] _pointer_data_40;
  assign _pointer_data_40 = _times_data_39[7'sd63];
  wire signed [2-1:0] _cond_data_52;
  assign _cond_data_52 = (_pointer_data_40)? -2'sd1 : 1'sd0;
  wire signed [65-1:0] _plus_data_53;
  assign _plus_data_53 = _times_data_39 + __delay_data_830__delay_829__delay_828__delay_827_sll_45;
  wire signed [65-1:0] _plus_data_54;
  assign _plus_data_54 = _plus_data_53 + _cond_data_52;
  wire signed [64-1:0] _sra_data_55;
  assign _sra_data_55 = _plus_data_54 >>> __delay_data_834__delay_833__delay_832__delay_831__variable_38;
  reg signed [64-1:0] _cond_data_58;
  reg [1-1:0] _greaterthan_data_59;
  reg [1-1:0] _lessthan_data_63;
  reg [1-1:0] _greatereq_data_67;
  reg signed [64-1:0] __delay_data_839_cond_58;
  reg signed [64-1:0] _cond_data_61;
  reg signed [64-1:0] _cond_data_65;
  reg [1-1:0] __delay_data_840_greatereq_67;
  reg signed [32-1:0] _cond_data_69;
  wire signed [32-1:0] mul_rshift_round_clip_2_z_data;
  assign mul_rshift_round_clip_2_z_data = _cond_data_69;
  reg [33-1:0] _stream_conv2d_2_sink_50_sink_count;
  reg [5-1:0] _stream_conv2d_2_sink_50_sink_mode;
  reg [16-1:0] _stream_conv2d_2_sink_50_sink_generator_id;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_offset;
  reg [33-1:0] _stream_conv2d_2_sink_50_sink_size;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_stride;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_2_sink_50_sink_size_buf;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_2_sink_50_sink_sel;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_waddr;
  reg _stream_conv2d_2_sink_50_sink_wenable;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_wdata;
  reg _stream_conv2d_2_sink_50_sink_fifo_enq;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_fifo_wdata;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_immediate;
  reg [33-1:0] _stream_conv2d_2_sink_51_sink_count;
  reg [5-1:0] _stream_conv2d_2_sink_51_sink_mode;
  reg [16-1:0] _stream_conv2d_2_sink_51_sink_generator_id;
  reg [32-1:0] _stream_conv2d_2_sink_51_sink_offset;
  reg [33-1:0] _stream_conv2d_2_sink_51_sink_size;
  reg [32-1:0] _stream_conv2d_2_sink_51_sink_stride;
  reg [32-1:0] _stream_conv2d_2_sink_51_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_2_sink_51_sink_size_buf;
  reg [32-1:0] _stream_conv2d_2_sink_51_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_2_sink_51_sink_sel;
  reg [32-1:0] _stream_conv2d_2_sink_51_sink_waddr;
  reg _stream_conv2d_2_sink_51_sink_wenable;
  reg [1-1:0] _stream_conv2d_2_sink_51_sink_wdata;
  reg _stream_conv2d_2_sink_51_sink_fifo_enq;
  reg [1-1:0] _stream_conv2d_2_sink_51_sink_fifo_wdata;
  reg [1-1:0] _stream_conv2d_2_sink_51_sink_immediate;
  reg _stream_celu_3_stream_ivalid;
  wire _stream_celu_3_stream_oready;
  wire _stream_celu_3_stream_internal_oready;
  assign _stream_celu_3_stream_internal_oready = 1;
  assign _stream_celu_3_stream_oready = _stream_celu_3_stream_internal_oready;
  reg [32-1:0] _stream_celu_3_fsm;
  localparam _stream_celu_3_fsm_init = 0;
  wire _stream_celu_3_run_flag;
  reg _stream_celu_3_source_start;
  wire _stream_celu_3_source_stop;
  reg _stream_celu_3_source_busy;
  wire _stream_celu_3_sink_start;
  wire _stream_celu_3_sink_stop;
  wire _stream_celu_3_sink_busy;
  wire _stream_celu_3_busy;
  reg _stream_celu_3_busy_reg;
  wire _stream_celu_3_is_root;
  assign _stream_celu_3_is_root = 1;
  reg [1-1:0] _stream_celu_3_parameter_0_next_parameter_data;
  reg _stream_celu_3_source_1_idle;
  reg [33-1:0] _stream_celu_3_source_1_source_count;
  reg [5-1:0] _stream_celu_3_source_1_source_mode;
  reg [16-1:0] _stream_celu_3_source_1_source_generator_id;
  reg [32-1:0] _stream_celu_3_source_1_source_offset;
  reg [33-1:0] _stream_celu_3_source_1_source_size;
  reg [32-1:0] _stream_celu_3_source_1_source_stride;
  reg [32-1:0] _stream_celu_3_source_1_source_offset_buf;
  reg [33-1:0] _stream_celu_3_source_1_source_size_buf;
  reg [32-1:0] _stream_celu_3_source_1_source_stride_buf;
  reg [8-1:0] _stream_celu_3_source_1_source_sel;
  reg [32-1:0] _stream_celu_3_source_1_source_ram_raddr;
  reg _stream_celu_3_source_1_source_ram_renable;
  wire [32-1:0] _stream_celu_3_source_1_source_ram_rdata;
  reg _stream_celu_3_source_1_source_fifo_deq;
  wire [32-1:0] _stream_celu_3_source_1_source_fifo_rdata;
  reg [32-1:0] _stream_celu_3_source_1_source_empty_data;
  reg [33-1:0] _stream_celu_3_sink_2_sink_count;
  reg [5-1:0] _stream_celu_3_sink_2_sink_mode;
  reg [16-1:0] _stream_celu_3_sink_2_sink_generator_id;
  reg [32-1:0] _stream_celu_3_sink_2_sink_offset;
  reg [33-1:0] _stream_celu_3_sink_2_sink_size;
  reg [32-1:0] _stream_celu_3_sink_2_sink_stride;
  reg [32-1:0] _stream_celu_3_sink_2_sink_offset_buf;
  reg [33-1:0] _stream_celu_3_sink_2_sink_size_buf;
  reg [32-1:0] _stream_celu_3_sink_2_sink_stride_buf;
  reg [8-1:0] _stream_celu_3_sink_2_sink_sel;
  reg [32-1:0] _stream_celu_3_sink_2_sink_waddr;
  reg _stream_celu_3_sink_2_sink_wenable;
  reg [32-1:0] _stream_celu_3_sink_2_sink_wdata;
  reg _stream_celu_3_sink_2_sink_fifo_enq;
  reg [32-1:0] _stream_celu_3_sink_2_sink_fifo_wdata;
  reg [32-1:0] _stream_celu_3_sink_2_sink_immediate;
  reg [32-1:0] main_fsm;
  localparam main_fsm_init = 0;
  reg [32-1:0] internal_state_counter;
  reg [32-1:0] conv2d_2_objaddr;
  reg [32-1:0] conv2d_2_arg_objaddr_0;
  reg [32-1:0] conv2d_2_arg_objaddr_1;
  reg [32-1:0] control_conv2d_2;
  localparam control_conv2d_2_init = 0;
  reg _control_conv2d_2_called;
  wire signed [32-1:0] conv2d_2_act_base_offset;
  reg signed [32-1:0] conv2d_2_act_base_offset_row;
  reg signed [32-1:0] conv2d_2_act_base_offset_bat;
  assign conv2d_2_act_base_offset = conv2d_2_act_base_offset_row + conv2d_2_act_base_offset_bat;
  reg signed [32-1:0] conv2d_2_filter_base_offset;
  reg [32-1:0] conv2d_2_next_stream_num_ops;
  wire signed [32-1:0] conv2d_2_out_base_offset;
  reg signed [32-1:0] conv2d_2_out_base_offset_val;
  reg signed [32-1:0] conv2d_2_out_base_offset_col;
  reg signed [32-1:0] conv2d_2_out_base_offset_row;
  reg signed [32-1:0] conv2d_2_out_base_offset_bat;
  reg signed [32-1:0] conv2d_2_out_base_offset_och;
  assign conv2d_2_out_base_offset = conv2d_2_out_base_offset_val + conv2d_2_out_base_offset_col + conv2d_2_out_base_offset_row + conv2d_2_out_base_offset_bat + conv2d_2_out_base_offset_och;
  reg conv2d_2_dma_flag_0;
  reg conv2d_2_dma_flag_1;
  reg conv2d_2_dma_flag_2;
  reg [32-1:0] conv2d_2_sync_comp_count;
  reg [32-1:0] conv2d_2_sync_out_count;
  reg [32-1:0] conv2d_2_write_count;
  reg [32-1:0] conv2d_2_next_out_write_size;
  reg [32-1:0] conv2d_2_col_count;
  reg [32-1:0] conv2d_2_row_count;
  reg [32-1:0] conv2d_2_bat_count;
  reg [32-1:0] conv2d_2_och_count;
  reg [2-1:0] conv2d_2_col_select;
  reg [2-1:0] conv2d_2_row_select;
  reg [32-1:0] conv2d_2_out_col_count;
  reg [32-1:0] conv2d_2_out_row_count;
  reg [32-1:0] conv2d_2_out_ram_select;
  reg [32-1:0] conv2d_2_prev_col_count;
  reg [32-1:0] conv2d_2_prev_row_count;
  reg [32-1:0] conv2d_2_prev_bat_count;
  reg [32-1:0] conv2d_2_prev_och_count;
  reg [2-1:0] conv2d_2_prev_row_select;
  reg [32-1:0] conv2d_2_stream_act_local_0;
  reg [32-1:0] conv2d_2_stream_act_local_1;
  reg [32-1:0] conv2d_2_stream_act_local_2;
  reg [32-1:0] conv2d_2_stream_act_local_3;
  reg [32-1:0] conv2d_2_stream_act_local_4;
  reg [32-1:0] conv2d_2_stream_act_local_5;
  reg [32-1:0] conv2d_2_stream_act_local_6;
  reg [32-1:0] conv2d_2_stream_act_local_7;
  reg [32-1:0] conv2d_2_stream_act_local_8;
  reg [32-1:0] conv2d_2_stream_out_local_val;
  reg [32-1:0] conv2d_2_stream_out_local_col;
  wire [32-1:0] conv2d_2_stream_out_local;
  assign conv2d_2_stream_out_local = conv2d_2_stream_out_local_val + conv2d_2_stream_out_local_col;
  reg [32-1:0] conv2d_2_act_page_comp_offset_0;
  reg [32-1:0] conv2d_2_act_page_comp_offset_1;
  reg [32-1:0] conv2d_2_act_page_comp_offset_2;
  reg [32-1:0] conv2d_2_act_page_dma_offset_0;
  reg [32-1:0] conv2d_2_act_page_dma_offset_1;
  reg [32-1:0] conv2d_2_act_page_dma_offset_2;
  reg [32-1:0] conv2d_2_filter_page_comp_offset;
  reg [32-1:0] conv2d_2_filter_page_dma_offset;
  reg conv2d_2_out_page;
  reg [32-1:0] conv2d_2_out_page_comp_offset;
  reg [32-1:0] conv2d_2_out_page_dma_offset;
  reg [32-1:0] conv2d_2_out_laddr_offset;
  reg conv2d_2_skip_read_filter;
  reg conv2d_2_skip_read_act;
  reg conv2d_2_skip_comp;
  reg conv2d_2_skip_write_out;
  wire [32-1:0] mask_addr_shifted_25;
  assign mask_addr_shifted_25 = conv2d_2_arg_objaddr_1 + conv2d_2_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_26;
  assign mask_addr_masked_26 = mask_addr_shifted_25 << 2;
  reg [32-1:0] _maxi_read_req_fsm;
  localparam _maxi_read_req_fsm_init = 0;
  reg [33-1:0] _maxi_read_cur_global_size;
  reg _maxi_read_cont;
  wire [8-1:0] pack_read_req_op_sel_27;
  wire [32-1:0] pack_read_req_local_addr_28;
  wire [32-1:0] pack_read_req_local_stride_29;
  wire [33-1:0] pack_read_req_local_size_30;
  wire [32-1:0] pack_read_req_local_blocksize_31;
  assign pack_read_req_op_sel_27 = _maxi_read_op_sel;
  assign pack_read_req_local_addr_28 = _maxi_read_local_addr;
  assign pack_read_req_local_stride_29 = _maxi_read_local_stride;
  assign pack_read_req_local_size_30 = _maxi_read_local_size;
  assign pack_read_req_local_blocksize_31 = _maxi_read_local_blocksize;
  wire [137-1:0] pack_read_req_packed_32;
  assign pack_read_req_packed_32 = { pack_read_req_op_sel_27, pack_read_req_local_addr_28, pack_read_req_local_stride_29, pack_read_req_local_size_30, pack_read_req_local_blocksize_31 };
  assign _maxi_read_req_fifo_wdata = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? pack_read_req_packed_32 : 'hx;
  assign _maxi_read_req_fifo_enq = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? (_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full && !_maxi_read_req_fifo_almost_full : 0;
  localparam _tmp_33 = 1;
  wire [_tmp_33-1:0] _tmp_34;
  assign _tmp_34 = !_maxi_read_req_fifo_almost_full;
  reg [_tmp_33-1:0] __tmp_34_1;
  wire [32-1:0] mask_addr_shifted_35;
  assign mask_addr_shifted_35 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_36;
  assign mask_addr_masked_36 = mask_addr_shifted_35 << 2;
  wire [32-1:0] mask_addr_shifted_37;
  assign mask_addr_shifted_37 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_38;
  assign mask_addr_masked_38 = mask_addr_shifted_37 << 2;
  wire [32-1:0] mask_addr_shifted_39;
  assign mask_addr_shifted_39 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_40;
  assign mask_addr_masked_40 = mask_addr_shifted_39 << 2;
  wire [32-1:0] mask_addr_shifted_41;
  assign mask_addr_shifted_41 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_42;
  assign mask_addr_masked_42 = mask_addr_shifted_41 << 2;
  wire [32-1:0] mask_addr_shifted_43;
  assign mask_addr_shifted_43 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_44;
  assign mask_addr_masked_44 = mask_addr_shifted_43 << 2;
  wire [32-1:0] mask_addr_shifted_45;
  assign mask_addr_shifted_45 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_46;
  assign mask_addr_masked_46 = mask_addr_shifted_45 << 2;
  reg _maxi_cond_0_1;
  reg [32-1:0] _maxi_read_data_fsm;
  localparam _maxi_read_data_fsm_init = 0;
  wire write_burst_block_ram_wvalid_47;
  wire write_burst_block_ram_wquit_48;
  reg [32-1:0] write_burst_fsm_0;
  localparam write_burst_fsm_0_init = 0;
  reg [7-1:0] write_burst_addr_49;
  reg [7-1:0] write_burst_stride_50;
  reg [33-1:0] write_burst_length_51;
  reg write_burst_done_52;
  assign ram_w32_l128_id1_1_wdata = ((write_burst_fsm_0 == 1) && write_burst_block_ram_wvalid_47)? maxi_rdata : 'hx;
  assign ram_w32_l128_id1_1_wenable = ((write_burst_fsm_0 == 1) && write_burst_block_ram_wvalid_47)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_53;
  wire write_burst_block_ram_wquit_54;
  reg [32-1:0] write_burst_fsm_1;
  localparam write_burst_fsm_1_init = 0;
  reg [7-1:0] write_burst_addr_55;
  reg [7-1:0] write_burst_stride_56;
  reg [33-1:0] write_burst_length_57;
  reg write_burst_done_58;
  assign ram_w32_l128_id2_1_addr = ((write_burst_fsm_1 == 1) && write_burst_block_ram_wvalid_53)? write_burst_addr_55 : 'hx;
  assign ram_w32_l128_id2_1_wdata = ((write_burst_fsm_1 == 1) && write_burst_block_ram_wvalid_53)? maxi_rdata : 'hx;
  assign ram_w32_l128_id2_1_wenable = ((write_burst_fsm_1 == 1) && write_burst_block_ram_wvalid_53)? 1'd1 : 0;
  assign ram_w32_l128_id2_1_enable = ((write_burst_fsm_1 == 1) && write_burst_block_ram_wvalid_53)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_59;
  wire write_burst_block_ram_wquit_60;
  reg [32-1:0] write_burst_fsm_2;
  localparam write_burst_fsm_2_init = 0;
  reg [7-1:0] write_burst_addr_61;
  reg [7-1:0] write_burst_stride_62;
  reg [33-1:0] write_burst_length_63;
  reg write_burst_done_64;
  assign ram_w32_l128_id3_1_addr = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_59)? write_burst_addr_61 : 'hx;
  assign ram_w32_l128_id3_1_wdata = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_59)? maxi_rdata : 'hx;
  assign ram_w32_l128_id3_1_wenable = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_59)? 1'd1 : 0;
  assign ram_w32_l128_id3_1_enable = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_59)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_65;
  wire write_burst_block_ram_wquit_66;
  reg [32-1:0] write_burst_fsm_3;
  localparam write_burst_fsm_3_init = 0;
  reg [7-1:0] write_burst_addr_67;
  reg [7-1:0] write_burst_stride_68;
  reg [33-1:0] write_burst_length_69;
  reg write_burst_done_70;
  assign ram_w32_l128_id4_1_addr = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_65)? write_burst_addr_67 : 'hx;
  assign ram_w32_l128_id4_1_wdata = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_65)? maxi_rdata : 'hx;
  assign ram_w32_l128_id4_1_wenable = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_65)? 1'd1 : 0;
  assign ram_w32_l128_id4_1_enable = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_65)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_71;
  wire write_burst_block_ram_wquit_72;
  reg [32-1:0] write_burst_fsm_4;
  localparam write_burst_fsm_4_init = 0;
  reg [7-1:0] write_burst_addr_73;
  reg [7-1:0] write_burst_stride_74;
  reg [33-1:0] write_burst_length_75;
  reg write_burst_done_76;
  assign ram_w32_l128_id5_1_addr = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_71)? write_burst_addr_73 : 'hx;
  assign ram_w32_l128_id5_1_wdata = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_71)? maxi_rdata : 'hx;
  assign ram_w32_l128_id5_1_wenable = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_71)? 1'd1 : 0;
  assign ram_w32_l128_id5_1_enable = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_71)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_77;
  wire write_burst_block_ram_wquit_78;
  reg [32-1:0] write_burst_fsm_5;
  localparam write_burst_fsm_5_init = 0;
  reg [7-1:0] write_burst_addr_79;
  reg [7-1:0] write_burst_stride_80;
  reg [33-1:0] write_burst_length_81;
  reg write_burst_done_82;
  assign ram_w32_l128_id6_1_addr = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_77)? write_burst_addr_79 : 'hx;
  assign ram_w32_l128_id6_1_wdata = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_77)? maxi_rdata : 'hx;
  assign ram_w32_l128_id6_1_wenable = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_77)? 1'd1 : 0;
  assign ram_w32_l128_id6_1_enable = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_77)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_83;
  wire write_burst_block_ram_wquit_84;
  reg [32-1:0] write_burst_fsm_6;
  localparam write_burst_fsm_6_init = 0;
  reg [7-1:0] write_burst_addr_85;
  reg [7-1:0] write_burst_stride_86;
  reg [33-1:0] write_burst_length_87;
  reg write_burst_done_88;
  assign ram_w32_l128_id7_1_addr = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_83)? write_burst_addr_85 : 'hx;
  assign ram_w32_l128_id7_1_wdata = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_83)? maxi_rdata : 'hx;
  assign ram_w32_l128_id7_1_wenable = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_83)? 1'd1 : 0;
  assign ram_w32_l128_id7_1_enable = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_83)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_89;
  wire write_burst_block_ram_wquit_90;
  reg [32-1:0] write_burst_fsm_7;
  localparam write_burst_fsm_7_init = 0;
  reg [7-1:0] write_burst_addr_91;
  reg [7-1:0] write_burst_stride_92;
  reg [33-1:0] write_burst_length_93;
  reg write_burst_done_94;
  assign ram_w32_l128_id8_1_addr = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_89)? write_burst_addr_91 : 'hx;
  assign ram_w32_l128_id8_1_wdata = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_89)? maxi_rdata : 'hx;
  assign ram_w32_l128_id8_1_wenable = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_89)? 1'd1 : 0;
  assign ram_w32_l128_id8_1_enable = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_89)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_95;
  wire write_burst_block_ram_wquit_96;
  reg [32-1:0] write_burst_fsm_8;
  localparam write_burst_fsm_8_init = 0;
  reg [7-1:0] write_burst_addr_97;
  reg [7-1:0] write_burst_stride_98;
  reg [33-1:0] write_burst_length_99;
  reg write_burst_done_100;
  assign ram_w32_l128_id9_1_addr = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_95)? write_burst_addr_97 : 'hx;
  assign ram_w32_l128_id9_1_wdata = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_95)? maxi_rdata : 'hx;
  assign ram_w32_l128_id9_1_wenable = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_95)? 1'd1 : 0;
  assign ram_w32_l128_id9_1_enable = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_95)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_9;
  localparam write_burst_block_fsm_9_init = 0;
  reg [33-1:0] write_burst_block_length_101;
  reg [32-1:0] write_burst_block_blocksize_102;
  reg write_burst_block_done_103;
  reg [32-1:0] write_burst_block_count_104;
  assign write_burst_block_ram_wvalid_47 = maxi_rvalid && (write_burst_block_fsm_9 == 1);
  assign write_burst_block_ram_wquit_48 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_53 = maxi_rvalid && (write_burst_block_fsm_9 == 2);
  assign write_burst_block_ram_wquit_54 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_59 = maxi_rvalid && (write_burst_block_fsm_9 == 3);
  assign write_burst_block_ram_wquit_60 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_65 = maxi_rvalid && (write_burst_block_fsm_9 == 4);
  assign write_burst_block_ram_wquit_66 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_71 = maxi_rvalid && (write_burst_block_fsm_9 == 5);
  assign write_burst_block_ram_wquit_72 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_77 = maxi_rvalid && (write_burst_block_fsm_9 == 6);
  assign write_burst_block_ram_wquit_78 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_83 = maxi_rvalid && (write_burst_block_fsm_9 == 7);
  assign write_burst_block_ram_wquit_84 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_89 = maxi_rvalid && (write_burst_block_fsm_9 == 8);
  assign write_burst_block_ram_wquit_90 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  assign write_burst_block_ram_wvalid_95 = maxi_rvalid && (write_burst_block_fsm_9 == 9);
  assign write_burst_block_ram_wquit_96 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_101 <= 1);
  wire [32-1:0] conv2d_2_mux_act_gaddr_0;
  assign conv2d_2_mux_act_gaddr_0 = (conv2d_2_row_select == 0)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_0) : 
                                    (conv2d_2_row_select == 1)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_2) : 
                                    (conv2d_2_row_select == 2)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_1) : 1'd0;
  wire [32-1:0] conv2d_2_mux_act_gaddr_1;
  assign conv2d_2_mux_act_gaddr_1 = (conv2d_2_row_select == 0)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_1) : 
                                    (conv2d_2_row_select == 1)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_0) : 
                                    (conv2d_2_row_select == 2)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_2) : 1'd0;
  wire [32-1:0] conv2d_2_mux_act_gaddr_2;
  assign conv2d_2_mux_act_gaddr_2 = (conv2d_2_row_select == 0)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_2) : 
                                    (conv2d_2_row_select == 1)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_1) : 
                                    (conv2d_2_row_select == 2)? conv2d_2_arg_objaddr_0 + (conv2d_2_act_base_offset + cparam_conv2d_2_act_offset_values_0) : 1'd0;
  wire conv2d_2_dma_pad_mask_0;
  assign conv2d_2_dma_pad_mask_0 = (conv2d_2_row_count + 0 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count + 0 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_dma_pad_mask_1;
  assign conv2d_2_dma_pad_mask_1 = (conv2d_2_row_count + 1 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count + 1 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_dma_pad_mask_2;
  assign conv2d_2_dma_pad_mask_2 = (conv2d_2_row_count + 2 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count + 2 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_mux_dma_pad_mask_0;
  assign conv2d_2_mux_dma_pad_mask_0 = (conv2d_2_row_select == 0)? conv2d_2_dma_pad_mask_0 : 
                                       (conv2d_2_row_select == 1)? conv2d_2_dma_pad_mask_2 : 
                                       (conv2d_2_row_select == 2)? conv2d_2_dma_pad_mask_1 : 1'd0;
  wire conv2d_2_mux_dma_pad_mask_1;
  assign conv2d_2_mux_dma_pad_mask_1 = (conv2d_2_row_select == 0)? conv2d_2_dma_pad_mask_1 : 
                                       (conv2d_2_row_select == 1)? conv2d_2_dma_pad_mask_0 : 
                                       (conv2d_2_row_select == 2)? conv2d_2_dma_pad_mask_2 : 1'd0;
  wire conv2d_2_mux_dma_pad_mask_2;
  assign conv2d_2_mux_dma_pad_mask_2 = (conv2d_2_row_select == 0)? conv2d_2_dma_pad_mask_2 : 
                                       (conv2d_2_row_select == 1)? conv2d_2_dma_pad_mask_1 : 
                                       (conv2d_2_row_select == 2)? conv2d_2_dma_pad_mask_0 : 1'd0;
  wire conv2d_2_mux_dma_flag_0;
  assign conv2d_2_mux_dma_flag_0 = (conv2d_2_prev_row_select == 0)? conv2d_2_dma_flag_0 : 
                                   (conv2d_2_prev_row_select == 1)? conv2d_2_dma_flag_2 : 
                                   (conv2d_2_prev_row_select == 2)? conv2d_2_dma_flag_1 : 1'd0;
  wire conv2d_2_mux_dma_flag_1;
  assign conv2d_2_mux_dma_flag_1 = (conv2d_2_prev_row_select == 0)? conv2d_2_dma_flag_1 : 
                                   (conv2d_2_prev_row_select == 1)? conv2d_2_dma_flag_0 : 
                                   (conv2d_2_prev_row_select == 2)? conv2d_2_dma_flag_2 : 1'd0;
  wire conv2d_2_mux_dma_flag_2;
  assign conv2d_2_mux_dma_flag_2 = (conv2d_2_prev_row_select == 0)? conv2d_2_dma_flag_2 : 
                                   (conv2d_2_prev_row_select == 1)? conv2d_2_dma_flag_1 : 
                                   (conv2d_2_prev_row_select == 2)? conv2d_2_dma_flag_0 : 1'd0;
  wire [32-1:0] mask_addr_shifted_105;
  assign mask_addr_shifted_105 = conv2d_2_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_106;
  assign mask_addr_masked_106 = mask_addr_shifted_105 << 2;
  wire write_burst_block_ram_wvalid_107;
  wire write_burst_block_ram_wquit_108;
  reg [32-1:0] write_burst_fsm_10;
  localparam write_burst_fsm_10_init = 0;
  reg [7-1:0] write_burst_addr_109;
  reg [7-1:0] write_burst_stride_110;
  reg [33-1:0] write_burst_length_111;
  reg write_burst_done_112;
  assign ram_w32_l128_id10_1_addr = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_107)? write_burst_addr_109 : 'hx;
  assign ram_w32_l128_id10_1_wdata = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_107)? maxi_rdata : 'hx;
  assign ram_w32_l128_id10_1_wenable = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_107)? 1'd1 : 0;
  assign ram_w32_l128_id10_1_enable = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_107)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_113;
  wire write_burst_block_ram_wquit_114;
  reg [32-1:0] write_burst_fsm_11;
  localparam write_burst_fsm_11_init = 0;
  reg [7-1:0] write_burst_addr_115;
  reg [7-1:0] write_burst_stride_116;
  reg [33-1:0] write_burst_length_117;
  reg write_burst_done_118;
  assign ram_w32_l128_id11_1_addr = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_113)? write_burst_addr_115 : 'hx;
  assign ram_w32_l128_id11_1_wdata = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_113)? maxi_rdata : 'hx;
  assign ram_w32_l128_id11_1_wenable = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_113)? 1'd1 : 0;
  assign ram_w32_l128_id11_1_enable = ((write_burst_fsm_11 == 1) && write_burst_block_ram_wvalid_113)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_119;
  wire write_burst_block_ram_wquit_120;
  reg [32-1:0] write_burst_fsm_12;
  localparam write_burst_fsm_12_init = 0;
  reg [7-1:0] write_burst_addr_121;
  reg [7-1:0] write_burst_stride_122;
  reg [33-1:0] write_burst_length_123;
  reg write_burst_done_124;
  assign ram_w32_l128_id12_1_addr = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_119)? write_burst_addr_121 : 'hx;
  assign ram_w32_l128_id12_1_wdata = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_119)? maxi_rdata : 'hx;
  assign ram_w32_l128_id12_1_wenable = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  assign ram_w32_l128_id12_1_enable = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_13;
  localparam write_burst_block_fsm_13_init = 0;
  reg [33-1:0] write_burst_block_length_125;
  reg [32-1:0] write_burst_block_blocksize_126;
  reg write_burst_block_done_127;
  reg [32-1:0] write_burst_block_count_128;
  assign write_burst_block_ram_wvalid_107 = maxi_rvalid && (write_burst_block_fsm_13 == 1);
  assign write_burst_block_ram_wquit_108 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_125 <= 1);
  assign write_burst_block_ram_wvalid_113 = maxi_rvalid && (write_burst_block_fsm_13 == 2);
  assign write_burst_block_ram_wquit_114 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_125 <= 1);
  assign write_burst_block_ram_wvalid_119 = maxi_rvalid && (write_burst_block_fsm_13 == 3);
  assign write_burst_block_ram_wquit_120 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_125 <= 1);
  wire [32-1:0] mask_addr_shifted_129;
  assign mask_addr_shifted_129 = conv2d_2_mux_act_gaddr_1 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_130;
  assign mask_addr_masked_130 = mask_addr_shifted_129 << 2;
  wire write_burst_block_ram_wvalid_131;
  wire write_burst_block_ram_wquit_132;
  reg [32-1:0] write_burst_fsm_14;
  localparam write_burst_fsm_14_init = 0;
  reg [7-1:0] write_burst_addr_133;
  reg [7-1:0] write_burst_stride_134;
  reg [33-1:0] write_burst_length_135;
  reg write_burst_done_136;
  assign ram_w32_l128_id13_1_addr = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_131)? write_burst_addr_133 : 'hx;
  assign ram_w32_l128_id13_1_wdata = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_131)? maxi_rdata : 'hx;
  assign ram_w32_l128_id13_1_wenable = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_131)? 1'd1 : 0;
  assign ram_w32_l128_id13_1_enable = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_131)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_137;
  wire write_burst_block_ram_wquit_138;
  reg [32-1:0] write_burst_fsm_15;
  localparam write_burst_fsm_15_init = 0;
  reg [7-1:0] write_burst_addr_139;
  reg [7-1:0] write_burst_stride_140;
  reg [33-1:0] write_burst_length_141;
  reg write_burst_done_142;
  assign ram_w32_l128_id14_1_addr = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_137)? write_burst_addr_139 : 'hx;
  assign ram_w32_l128_id14_1_wdata = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_137)? maxi_rdata : 'hx;
  assign ram_w32_l128_id14_1_wenable = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_137)? 1'd1 : 0;
  assign ram_w32_l128_id14_1_enable = ((write_burst_fsm_15 == 1) && write_burst_block_ram_wvalid_137)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_143;
  wire write_burst_block_ram_wquit_144;
  reg [32-1:0] write_burst_fsm_16;
  localparam write_burst_fsm_16_init = 0;
  reg [7-1:0] write_burst_addr_145;
  reg [7-1:0] write_burst_stride_146;
  reg [33-1:0] write_burst_length_147;
  reg write_burst_done_148;
  assign ram_w32_l128_id15_1_addr = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_143)? write_burst_addr_145 : 'hx;
  assign ram_w32_l128_id15_1_wdata = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_143)? maxi_rdata : 'hx;
  assign ram_w32_l128_id15_1_wenable = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_143)? 1'd1 : 0;
  assign ram_w32_l128_id15_1_enable = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_143)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_17;
  localparam write_burst_block_fsm_17_init = 0;
  reg [33-1:0] write_burst_block_length_149;
  reg [32-1:0] write_burst_block_blocksize_150;
  reg write_burst_block_done_151;
  reg [32-1:0] write_burst_block_count_152;
  assign write_burst_block_ram_wvalid_131 = maxi_rvalid && (write_burst_block_fsm_17 == 1);
  assign write_burst_block_ram_wquit_132 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_149 <= 1);
  assign write_burst_block_ram_wvalid_137 = maxi_rvalid && (write_burst_block_fsm_17 == 2);
  assign write_burst_block_ram_wquit_138 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_149 <= 1);
  assign write_burst_block_ram_wvalid_143 = maxi_rvalid && (write_burst_block_fsm_17 == 3);
  assign write_burst_block_ram_wquit_144 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_149 <= 1);
  wire [32-1:0] mask_addr_shifted_153;
  assign mask_addr_shifted_153 = conv2d_2_mux_act_gaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_154;
  assign mask_addr_masked_154 = mask_addr_shifted_153 << 2;
  wire write_burst_block_ram_wvalid_155;
  wire write_burst_block_ram_wquit_156;
  reg [32-1:0] write_burst_fsm_18;
  localparam write_burst_fsm_18_init = 0;
  reg [7-1:0] write_burst_addr_157;
  reg [7-1:0] write_burst_stride_158;
  reg [33-1:0] write_burst_length_159;
  reg write_burst_done_160;
  assign ram_w32_l128_id16_1_addr = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_155)? write_burst_addr_157 : 'hx;
  assign ram_w32_l128_id16_1_wdata = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_155)? maxi_rdata : 'hx;
  assign ram_w32_l128_id16_1_wenable = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_155)? 1'd1 : 0;
  assign ram_w32_l128_id16_1_enable = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_155)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_161;
  wire write_burst_block_ram_wquit_162;
  reg [32-1:0] write_burst_fsm_19;
  localparam write_burst_fsm_19_init = 0;
  reg [7-1:0] write_burst_addr_163;
  reg [7-1:0] write_burst_stride_164;
  reg [33-1:0] write_burst_length_165;
  reg write_burst_done_166;
  assign ram_w32_l128_id17_1_addr = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_161)? write_burst_addr_163 : 'hx;
  assign ram_w32_l128_id17_1_wdata = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_161)? maxi_rdata : 'hx;
  assign ram_w32_l128_id17_1_wenable = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  assign ram_w32_l128_id17_1_enable = ((write_burst_fsm_19 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_167;
  wire write_burst_block_ram_wquit_168;
  reg [32-1:0] write_burst_fsm_20;
  localparam write_burst_fsm_20_init = 0;
  reg [7-1:0] write_burst_addr_169;
  reg [7-1:0] write_burst_stride_170;
  reg [33-1:0] write_burst_length_171;
  reg write_burst_done_172;
  assign ram_w32_l128_id18_1_addr = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_167)? write_burst_addr_169 : 'hx;
  assign ram_w32_l128_id18_1_wdata = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_167)? maxi_rdata : 'hx;
  assign ram_w32_l128_id18_1_wenable = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_167)? 1'd1 : 0;
  assign ram_w32_l128_id18_1_enable = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_167)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_21;
  localparam write_burst_block_fsm_21_init = 0;
  reg [33-1:0] write_burst_block_length_173;
  reg [32-1:0] write_burst_block_blocksize_174;
  reg write_burst_block_done_175;
  reg [32-1:0] write_burst_block_count_176;
  assign write_burst_block_ram_wvalid_155 = maxi_rvalid && (write_burst_block_fsm_21 == 1);
  assign write_burst_block_ram_wquit_156 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_173 <= 1);
  assign write_burst_block_ram_wvalid_161 = maxi_rvalid && (write_burst_block_fsm_21 == 2);
  assign write_burst_block_ram_wquit_162 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_173 <= 1);
  assign write_burst_block_ram_wvalid_167 = maxi_rvalid && (write_burst_block_fsm_21 == 3);
  assign write_burst_block_ram_wquit_168 = 0 || maxi_rvalid && 0 || maxi_rvalid && (write_burst_block_length_173 <= 1);
  reg [32-1:0] conv2d_2_comp_fsm;
  localparam conv2d_2_comp_fsm_init = 0;
  reg [32-1:0] conv2d_2_filter_page_comp_offset_buf;
  reg [32-1:0] conv2d_2_act_page_comp_offset_buf_0;
  reg [32-1:0] conv2d_2_act_page_comp_offset_buf_1;
  reg [32-1:0] conv2d_2_act_page_comp_offset_buf_2;
  reg [32-1:0] conv2d_2_out_page_comp_offset_buf;
  reg [32-1:0] conv2d_2_row_count_buf;
  reg [2-1:0] conv2d_2_row_select_buf;
  reg [32-1:0] conv2d_2_och_count_buf;
  wire conv2d_2_stream_pad_mask_0_0;
  assign conv2d_2_stream_pad_mask_0_0 = (conv2d_2_col_count + 0 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 0 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 0 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 0 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_0_1;
  assign conv2d_2_stream_pad_mask_0_1 = (conv2d_2_col_count + 1 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 1 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 0 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 0 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_0_2;
  assign conv2d_2_stream_pad_mask_0_2 = (conv2d_2_col_count + 2 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 2 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 0 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 0 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_1_0;
  assign conv2d_2_stream_pad_mask_1_0 = (conv2d_2_col_count + 0 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 0 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 1 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 1 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_1_1;
  assign conv2d_2_stream_pad_mask_1_1 = (conv2d_2_col_count + 1 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 1 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 1 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 1 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_1_2;
  assign conv2d_2_stream_pad_mask_1_2 = (conv2d_2_col_count + 2 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 2 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 1 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 1 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_2_0;
  assign conv2d_2_stream_pad_mask_2_0 = (conv2d_2_col_count + 0 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 0 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 2 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 2 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_2_1;
  assign conv2d_2_stream_pad_mask_2_1 = (conv2d_2_col_count + 1 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 1 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 2 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 2 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  wire conv2d_2_stream_pad_mask_2_2;
  assign conv2d_2_stream_pad_mask_2_2 = (conv2d_2_col_count + 2 < cparam_conv2d_2_pad_col_left) || (conv2d_2_col_count + 2 >= cparam_conv2d_2_act_num_col + cparam_conv2d_2_pad_col_left) || (conv2d_2_row_count_buf + 2 < cparam_conv2d_2_pad_row_top) || (conv2d_2_row_count_buf + 2 >= cparam_conv2d_2_act_num_row + cparam_conv2d_2_pad_row_top);
  reg [9-1:0] conv2d_2_stream_pad_masks;
  wire [4-1:0] stream_conv2d_2_parameter_0_data;
  wire [2-1:0] stream_conv2d_2_parameter_1_data;
  wire [2-1:0] stream_conv2d_2_parameter_2_data;
  wire [9-1:0] stream_conv2d_2_parameter_3_data;
  wire [1-1:0] stream_conv2d_2_parameter_4_data;
  wire [1-1:0] stream_conv2d_2__reduce_reset_data;
  wire [1-1:0] stream_conv2d_2_parameter_6_data;
  wire [32-1:0] stream_conv2d_2_source_7_data;
  wire [1-1:0] stream_conv2d_2_parameter_8_data;
  wire [32-1:0] stream_conv2d_2_source_9_data;
  wire [1-1:0] stream_conv2d_2_parameter_10_data;
  wire [32-1:0] stream_conv2d_2_source_11_data;
  wire [1-1:0] stream_conv2d_2_parameter_12_data;
  wire [32-1:0] stream_conv2d_2_source_13_data;
  wire [1-1:0] stream_conv2d_2_parameter_14_data;
  wire [32-1:0] stream_conv2d_2_source_15_data;
  wire [1-1:0] stream_conv2d_2_parameter_16_data;
  wire [1-1:0] stream_conv2d_2_parameter_17_data;
  wire [1-1:0] stream_conv2d_2_parameter_18_data;
  wire [1-1:0] stream_conv2d_2_parameter_19_data;
  wire [32-1:0] stream_conv2d_2_source_20_data;
  wire [32-1:0] stream_conv2d_2_source_21_data;
  wire [32-1:0] stream_conv2d_2_source_22_data;
  wire [32-1:0] stream_conv2d_2_source_23_data;
  wire [32-1:0] stream_conv2d_2_source_24_data;
  wire [32-1:0] stream_conv2d_2_source_25_data;
  wire [32-1:0] stream_conv2d_2_source_26_data;
  wire [32-1:0] stream_conv2d_2_source_27_data;
  wire [32-1:0] stream_conv2d_2_source_28_data;
  wire [32-1:0] stream_conv2d_2_source_29_data;
  wire [32-1:0] stream_conv2d_2_source_30_data;
  wire [32-1:0] stream_conv2d_2_source_31_data;
  wire [32-1:0] stream_conv2d_2_source_32_data;
  wire [32-1:0] stream_conv2d_2_source_33_data;
  wire [32-1:0] stream_conv2d_2_source_34_data;
  wire [32-1:0] stream_conv2d_2_source_35_data;
  wire [32-1:0] stream_conv2d_2_source_36_data;
  wire [32-1:0] stream_conv2d_2_source_37_data;
  reg __stream_conv2d_2_stream_ivalid_1;
  reg __stream_conv2d_2_stream_ivalid_2;
  reg __stream_conv2d_2_stream_ivalid_3;
  reg __stream_conv2d_2_stream_ivalid_4;
  reg __stream_conv2d_2_stream_ivalid_5;
  reg __stream_conv2d_2_stream_ivalid_6;
  reg __stream_conv2d_2_stream_ivalid_7;
  reg __stream_conv2d_2_stream_ivalid_8;
  reg __stream_conv2d_2_stream_ivalid_9;
  reg __stream_conv2d_2_stream_ivalid_10;
  reg __stream_conv2d_2_stream_ivalid_11;
  reg __stream_conv2d_2_stream_ivalid_12;
  reg __stream_conv2d_2_stream_ivalid_13;
  reg __stream_conv2d_2_stream_ivalid_14;
  reg __stream_conv2d_2_stream_ivalid_15;
  reg __stream_conv2d_2_stream_ivalid_16;
  reg __stream_conv2d_2_stream_ivalid_17;
  reg __stream_conv2d_2_stream_ivalid_18;
  reg __stream_conv2d_2_stream_ivalid_19;
  reg __stream_conv2d_2_stream_ivalid_20;
  reg __stream_conv2d_2_stream_ivalid_21;
  reg __stream_conv2d_2_stream_ivalid_22;
  reg __stream_conv2d_2_stream_ivalid_23;
  reg __stream_conv2d_2_stream_ivalid_24;
  reg __stream_conv2d_2_stream_ivalid_25;
  reg __stream_conv2d_2_stream_ivalid_26;
  reg __stream_conv2d_2_stream_ivalid_27;
  reg __stream_conv2d_2_stream_ivalid_28;
  reg __stream_conv2d_2_stream_ivalid_29;
  wire [32-1:0] _slice_data_278;
  assign _slice_data_278 = stream_conv2d_2_source_7_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_279;
  assign _reinterpretcast_src_279 = _slice_data_278;
  wire signed [32-1:0] _reinterpretcast_data_279;
  assign _reinterpretcast_data_279 = _reinterpretcast_src_279;
  wire signed [32-1:0] _cond_data_280;
  assign _cond_data_280 = (stream_conv2d_2_parameter_6_data)? _reinterpretcast_data_279 : _reinterpretcast_data_279;
  wire [32-1:0] _slice_data_285;
  assign _slice_data_285 = stream_conv2d_2_source_9_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_286;
  assign _reinterpretcast_src_286 = _slice_data_285;
  wire signed [32-1:0] _reinterpretcast_data_286;
  assign _reinterpretcast_data_286 = _reinterpretcast_src_286;
  wire signed [32-1:0] _cond_data_287;
  assign _cond_data_287 = (stream_conv2d_2_parameter_8_data)? _reinterpretcast_data_286 : _reinterpretcast_data_286;
  wire [32-1:0] _slice_data_292;
  assign _slice_data_292 = stream_conv2d_2_source_11_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_293;
  assign _reinterpretcast_src_293 = _slice_data_292;
  wire [32-1:0] _reinterpretcast_data_293;
  assign _reinterpretcast_data_293 = _reinterpretcast_src_293;
  wire [32-1:0] _cond_data_294;
  assign _cond_data_294 = (stream_conv2d_2_parameter_10_data)? _reinterpretcast_data_293 : _reinterpretcast_data_293;
  wire [32-1:0] _slice_data_299;
  assign _slice_data_299 = stream_conv2d_2_source_13_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_300;
  assign _reinterpretcast_src_300 = _slice_data_299;
  wire [32-1:0] _reinterpretcast_data_300;
  assign _reinterpretcast_data_300 = _reinterpretcast_src_300;
  wire [32-1:0] _cond_data_301;
  assign _cond_data_301 = (stream_conv2d_2_parameter_12_data)? _reinterpretcast_data_300 : _reinterpretcast_data_300;
  wire [32-1:0] _slice_data_306;
  assign _slice_data_306 = stream_conv2d_2_source_15_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_307;
  assign _reinterpretcast_src_307 = _slice_data_306;
  wire [32-1:0] _reinterpretcast_data_307;
  assign _reinterpretcast_data_307 = _reinterpretcast_src_307;
  wire [32-1:0] _cond_data_308;
  assign _cond_data_308 = (stream_conv2d_2_parameter_14_data)? _reinterpretcast_data_307 : _reinterpretcast_data_307;
  reg [1-1:0] _eq_data_322;
  reg [1-1:0] _eq_data_326;
  reg [1-1:0] _eq_data_329;
  reg [1-1:0] _eq_data_332;
  reg [1-1:0] _eq_data_336;
  reg [1-1:0] _eq_data_339;
  reg [1-1:0] _eq_data_342;
  reg [1-1:0] _eq_data_346;
  reg [1-1:0] _eq_data_349;
  reg [1-1:0] _eq_data_352;
  reg [1-1:0] _eq_data_356;
  reg [1-1:0] _eq_data_359;
  reg [1-1:0] _eq_data_362;
  reg [1-1:0] _eq_data_366;
  reg [1-1:0] _eq_data_369;
  reg [1-1:0] _eq_data_372;
  reg [1-1:0] _eq_data_376;
  reg [1-1:0] _eq_data_379;
  reg [1-1:0] _eq_data_382;
  reg [1-1:0] _eq_data_386;
  reg [1-1:0] _eq_data_389;
  reg [1-1:0] _eq_data_392;
  reg [1-1:0] _eq_data_396;
  reg [1-1:0] _eq_data_399;
  reg [1-1:0] _eq_data_402;
  reg [1-1:0] _eq_data_406;
  reg [1-1:0] _eq_data_409;
  reg [1-1:0] _eq_data_412;
  reg [1-1:0] _eq_data_416;
  reg [1-1:0] _eq_data_419;
  reg [1-1:0] _eq_data_422;
  reg [1-1:0] _eq_data_426;
  reg [1-1:0] _eq_data_429;
  reg [1-1:0] _eq_data_432;
  reg [1-1:0] _eq_data_436;
  reg [1-1:0] _eq_data_439;
  reg [1-1:0] _eq_data_442;
  reg [1-1:0] _eq_data_446;
  reg [1-1:0] _eq_data_449;
  reg [1-1:0] _eq_data_452;
  reg [1-1:0] _eq_data_456;
  reg [1-1:0] _eq_data_459;
  reg [1-1:0] _eq_data_462;
  reg [1-1:0] _eq_data_466;
  reg [1-1:0] _eq_data_469;
  reg [1-1:0] _eq_data_472;
  reg [1-1:0] _eq_data_476;
  reg [1-1:0] _eq_data_479;
  reg [1-1:0] _eq_data_482;
  reg [1-1:0] _eq_data_486;
  reg [1-1:0] _eq_data_489;
  reg [1-1:0] _eq_data_492;
  reg [1-1:0] _eq_data_496;
  reg [1-1:0] _eq_data_499;
  wire [32-1:0] _reinterpretcast_src_592;
  assign _reinterpretcast_src_592 = stream_conv2d_2_source_29_data;
  wire signed [32-1:0] _reinterpretcast_data_592;
  assign _reinterpretcast_data_592 = _reinterpretcast_src_592;
  wire [32-1:0] _reinterpretcast_src_593;
  assign _reinterpretcast_src_593 = stream_conv2d_2_source_30_data;
  wire signed [32-1:0] _reinterpretcast_data_593;
  assign _reinterpretcast_data_593 = _reinterpretcast_src_593;
  wire [32-1:0] _reinterpretcast_src_594;
  assign _reinterpretcast_src_594 = stream_conv2d_2_source_31_data;
  wire signed [32-1:0] _reinterpretcast_data_594;
  assign _reinterpretcast_data_594 = _reinterpretcast_src_594;
  wire [32-1:0] _reinterpretcast_src_595;
  assign _reinterpretcast_src_595 = stream_conv2d_2_source_32_data;
  wire signed [32-1:0] _reinterpretcast_data_595;
  assign _reinterpretcast_data_595 = _reinterpretcast_src_595;
  wire [32-1:0] _reinterpretcast_src_596;
  assign _reinterpretcast_src_596 = stream_conv2d_2_source_33_data;
  wire signed [32-1:0] _reinterpretcast_data_596;
  assign _reinterpretcast_data_596 = _reinterpretcast_src_596;
  wire [32-1:0] _reinterpretcast_src_597;
  assign _reinterpretcast_src_597 = stream_conv2d_2_source_34_data;
  wire signed [32-1:0] _reinterpretcast_data_597;
  assign _reinterpretcast_data_597 = _reinterpretcast_src_597;
  wire [32-1:0] _reinterpretcast_src_598;
  assign _reinterpretcast_src_598 = stream_conv2d_2_source_35_data;
  wire signed [32-1:0] _reinterpretcast_data_598;
  assign _reinterpretcast_data_598 = _reinterpretcast_src_598;
  wire [32-1:0] _reinterpretcast_src_599;
  assign _reinterpretcast_src_599 = stream_conv2d_2_source_36_data;
  wire signed [32-1:0] _reinterpretcast_data_599;
  assign _reinterpretcast_data_599 = _reinterpretcast_src_599;
  wire [32-1:0] _reinterpretcast_src_600;
  assign _reinterpretcast_src_600 = stream_conv2d_2_source_37_data;
  wire signed [32-1:0] _reinterpretcast_data_600;
  assign _reinterpretcast_data_600 = _reinterpretcast_src_600;
  wire [1-1:0] _pointer_data_601;
  assign _pointer_data_601 = stream_conv2d_2_parameter_3_data[1'sd0];
  wire [1-1:0] _pointer_data_603;
  assign _pointer_data_603 = stream_conv2d_2_parameter_3_data[2'sd1];
  wire [1-1:0] _pointer_data_605;
  assign _pointer_data_605 = stream_conv2d_2_parameter_3_data[3'sd2];
  wire [1-1:0] _pointer_data_607;
  assign _pointer_data_607 = stream_conv2d_2_parameter_3_data[3'sd3];
  wire [1-1:0] _pointer_data_609;
  assign _pointer_data_609 = stream_conv2d_2_parameter_3_data[4'sd4];
  wire [1-1:0] _pointer_data_611;
  assign _pointer_data_611 = stream_conv2d_2_parameter_3_data[4'sd5];
  wire [1-1:0] _pointer_data_613;
  assign _pointer_data_613 = stream_conv2d_2_parameter_3_data[4'sd6];
  wire [1-1:0] _pointer_data_615;
  assign _pointer_data_615 = stream_conv2d_2_parameter_3_data[4'sd7];
  wire [1-1:0] _pointer_data_617;
  assign _pointer_data_617 = stream_conv2d_2_parameter_3_data[5'sd8];
  reg [32-1:0] _plus_data_654;
  reg [32-1:0] _plus_data_673;
  reg [32-1:0] _plus_data_692;
  reg [32-1:0] _plus_data_711;
  reg [32-1:0] _plus_data_730;
  reg [32-1:0] _plus_data_749;
  reg [32-1:0] _plus_data_768;
  reg [32-1:0] _plus_data_787;
  reg [32-1:0] _plus_data_806;
  reg [32-1:0] _plus_data_822;
  reg [32-1:0] _plus_data_841;
  reg [32-1:0] __delay_data_866__variable_315;
  reg [32-1:0] __delay_data_867__variable_314;
  reg [32-1:0] __delay_data_868__variable_313;
  reg [32-1:0] __delay_data_869__variable_318;
  reg [32-1:0] __delay_data_870__variable_317;
  reg [32-1:0] __delay_data_871__variable_316;
  reg [32-1:0] __delay_data_872__variable_321;
  reg [32-1:0] __delay_data_873__variable_320;
  reg [32-1:0] __delay_data_874__variable_319;
  reg [1-1:0] __delay_data_875_pointer_601;
  reg signed [32-1:0] __delay_data_876_reinterpretcast_592;
  reg [1-1:0] __delay_data_877_pointer_603;
  reg signed [32-1:0] __delay_data_878_reinterpretcast_593;
  reg [1-1:0] __delay_data_879_pointer_605;
  reg signed [32-1:0] __delay_data_880_reinterpretcast_594;
  reg [1-1:0] __delay_data_881_pointer_607;
  reg signed [32-1:0] __delay_data_882_reinterpretcast_595;
  reg [1-1:0] __delay_data_883_pointer_609;
  reg signed [32-1:0] __delay_data_884_reinterpretcast_596;
  reg [1-1:0] __delay_data_885_pointer_611;
  reg signed [32-1:0] __delay_data_886_reinterpretcast_597;
  reg [1-1:0] __delay_data_887_pointer_613;
  reg signed [32-1:0] __delay_data_888_reinterpretcast_598;
  reg [1-1:0] __delay_data_889_pointer_615;
  reg signed [32-1:0] __delay_data_890_reinterpretcast_599;
  reg [1-1:0] __delay_data_891_pointer_617;
  reg signed [32-1:0] __delay_data_892_reinterpretcast_600;
  reg [1-1:0] __delay_data_893__variable_264;
  reg [4-1:0] __delay_data_918__variable_259;
  reg signed [32-1:0] __delay_data_931_cond_280;
  reg signed [32-1:0] __delay_data_950_cond_287;
  wire signed [32-1:0] _cond_data_324;
  assign _cond_data_324 = (_eq_data_322)? __delay_data_866__variable_315 : 1'sd0;
  wire signed [32-1:0] _cond_data_328;
  assign _cond_data_328 = (_eq_data_326)? __delay_data_867__variable_314 : _cond_data_324;
  wire signed [32-1:0] _cond_data_331;
  assign _cond_data_331 = (_eq_data_329)? __delay_data_868__variable_313 : _cond_data_328;
  wire signed [32-1:0] _cond_data_334;
  assign _cond_data_334 = (_eq_data_332)? __delay_data_868__variable_313 : 1'sd0;
  wire signed [32-1:0] _cond_data_338;
  assign _cond_data_338 = (_eq_data_336)? __delay_data_866__variable_315 : _cond_data_334;
  wire signed [32-1:0] _cond_data_341;
  assign _cond_data_341 = (_eq_data_339)? __delay_data_867__variable_314 : _cond_data_338;
  wire signed [32-1:0] _cond_data_344;
  assign _cond_data_344 = (_eq_data_342)? __delay_data_867__variable_314 : 1'sd0;
  wire signed [32-1:0] _cond_data_348;
  assign _cond_data_348 = (_eq_data_346)? __delay_data_868__variable_313 : _cond_data_344;
  wire signed [32-1:0] _cond_data_351;
  assign _cond_data_351 = (_eq_data_349)? __delay_data_866__variable_315 : _cond_data_348;
  wire signed [32-1:0] _cond_data_354;
  assign _cond_data_354 = (_eq_data_352)? __delay_data_869__variable_318 : 1'sd0;
  wire signed [32-1:0] _cond_data_358;
  assign _cond_data_358 = (_eq_data_356)? __delay_data_870__variable_317 : _cond_data_354;
  wire signed [32-1:0] _cond_data_361;
  assign _cond_data_361 = (_eq_data_359)? __delay_data_871__variable_316 : _cond_data_358;
  wire signed [32-1:0] _cond_data_364;
  assign _cond_data_364 = (_eq_data_362)? __delay_data_871__variable_316 : 1'sd0;
  wire signed [32-1:0] _cond_data_368;
  assign _cond_data_368 = (_eq_data_366)? __delay_data_869__variable_318 : _cond_data_364;
  wire signed [32-1:0] _cond_data_371;
  assign _cond_data_371 = (_eq_data_369)? __delay_data_870__variable_317 : _cond_data_368;
  wire signed [32-1:0] _cond_data_374;
  assign _cond_data_374 = (_eq_data_372)? __delay_data_870__variable_317 : 1'sd0;
  wire signed [32-1:0] _cond_data_378;
  assign _cond_data_378 = (_eq_data_376)? __delay_data_871__variable_316 : _cond_data_374;
  wire signed [32-1:0] _cond_data_381;
  assign _cond_data_381 = (_eq_data_379)? __delay_data_869__variable_318 : _cond_data_378;
  wire signed [32-1:0] _cond_data_384;
  assign _cond_data_384 = (_eq_data_382)? __delay_data_872__variable_321 : 1'sd0;
  wire signed [32-1:0] _cond_data_388;
  assign _cond_data_388 = (_eq_data_386)? __delay_data_873__variable_320 : _cond_data_384;
  wire signed [32-1:0] _cond_data_391;
  assign _cond_data_391 = (_eq_data_389)? __delay_data_874__variable_319 : _cond_data_388;
  wire signed [32-1:0] _cond_data_394;
  assign _cond_data_394 = (_eq_data_392)? __delay_data_874__variable_319 : 1'sd0;
  wire signed [32-1:0] _cond_data_398;
  assign _cond_data_398 = (_eq_data_396)? __delay_data_872__variable_321 : _cond_data_394;
  wire signed [32-1:0] _cond_data_401;
  assign _cond_data_401 = (_eq_data_399)? __delay_data_873__variable_320 : _cond_data_398;
  wire signed [32-1:0] _cond_data_404;
  assign _cond_data_404 = (_eq_data_402)? __delay_data_873__variable_320 : 1'sd0;
  wire signed [32-1:0] _cond_data_408;
  assign _cond_data_408 = (_eq_data_406)? __delay_data_874__variable_319 : _cond_data_404;
  wire signed [32-1:0] _cond_data_411;
  assign _cond_data_411 = (_eq_data_409)? __delay_data_872__variable_321 : _cond_data_408;
  wire signed [32-1:0] _cond_data_414;
  assign _cond_data_414 = (_eq_data_412)? _cond_data_391 : 1'sd0;
  wire signed [32-1:0] _cond_data_418;
  assign _cond_data_418 = (_eq_data_416)? _cond_data_361 : _cond_data_414;
  wire signed [32-1:0] _cond_data_421;
  assign _cond_data_421 = (_eq_data_419)? _cond_data_331 : _cond_data_418;
  wire signed [32-1:0] _cond_data_424;
  assign _cond_data_424 = (_eq_data_422)? _cond_data_331 : 1'sd0;
  wire signed [32-1:0] _cond_data_428;
  assign _cond_data_428 = (_eq_data_426)? _cond_data_391 : _cond_data_424;
  wire signed [32-1:0] _cond_data_431;
  assign _cond_data_431 = (_eq_data_429)? _cond_data_361 : _cond_data_428;
  wire signed [32-1:0] _cond_data_434;
  assign _cond_data_434 = (_eq_data_432)? _cond_data_361 : 1'sd0;
  wire signed [32-1:0] _cond_data_438;
  assign _cond_data_438 = (_eq_data_436)? _cond_data_331 : _cond_data_434;
  wire signed [32-1:0] _cond_data_441;
  assign _cond_data_441 = (_eq_data_439)? _cond_data_391 : _cond_data_438;
  wire signed [32-1:0] _cond_data_444;
  assign _cond_data_444 = (_eq_data_442)? _cond_data_401 : 1'sd0;
  wire signed [32-1:0] _cond_data_448;
  assign _cond_data_448 = (_eq_data_446)? _cond_data_371 : _cond_data_444;
  wire signed [32-1:0] _cond_data_451;
  assign _cond_data_451 = (_eq_data_449)? _cond_data_341 : _cond_data_448;
  wire signed [32-1:0] _cond_data_454;
  assign _cond_data_454 = (_eq_data_452)? _cond_data_341 : 1'sd0;
  wire signed [32-1:0] _cond_data_458;
  assign _cond_data_458 = (_eq_data_456)? _cond_data_401 : _cond_data_454;
  wire signed [32-1:0] _cond_data_461;
  assign _cond_data_461 = (_eq_data_459)? _cond_data_371 : _cond_data_458;
  wire signed [32-1:0] _cond_data_464;
  assign _cond_data_464 = (_eq_data_462)? _cond_data_371 : 1'sd0;
  wire signed [32-1:0] _cond_data_468;
  assign _cond_data_468 = (_eq_data_466)? _cond_data_341 : _cond_data_464;
  wire signed [32-1:0] _cond_data_471;
  assign _cond_data_471 = (_eq_data_469)? _cond_data_401 : _cond_data_468;
  wire signed [32-1:0] _cond_data_474;
  assign _cond_data_474 = (_eq_data_472)? _cond_data_411 : 1'sd0;
  wire signed [32-1:0] _cond_data_478;
  assign _cond_data_478 = (_eq_data_476)? _cond_data_381 : _cond_data_474;
  wire signed [32-1:0] _cond_data_481;
  assign _cond_data_481 = (_eq_data_479)? _cond_data_351 : _cond_data_478;
  wire signed [32-1:0] _cond_data_484;
  assign _cond_data_484 = (_eq_data_482)? _cond_data_351 : 1'sd0;
  wire signed [32-1:0] _cond_data_488;
  assign _cond_data_488 = (_eq_data_486)? _cond_data_411 : _cond_data_484;
  wire signed [32-1:0] _cond_data_491;
  assign _cond_data_491 = (_eq_data_489)? _cond_data_381 : _cond_data_488;
  wire signed [32-1:0] _cond_data_494;
  assign _cond_data_494 = (_eq_data_492)? _cond_data_381 : 1'sd0;
  wire signed [32-1:0] _cond_data_498;
  assign _cond_data_498 = (_eq_data_496)? _cond_data_351 : _cond_data_494;
  wire signed [32-1:0] _cond_data_501;
  assign _cond_data_501 = (_eq_data_499)? _cond_data_411 : _cond_data_498;
  wire signed [32-1:0] _reinterpretcast_src_538;
  assign _reinterpretcast_src_538 = _cond_data_421;
  wire signed [32-1:0] _reinterpretcast_data_538;
  assign _reinterpretcast_data_538 = _reinterpretcast_src_538;
  wire signed [32-1:0] _reinterpretcast_src_539;
  assign _reinterpretcast_src_539 = _cond_data_451;
  wire signed [32-1:0] _reinterpretcast_data_539;
  assign _reinterpretcast_data_539 = _reinterpretcast_src_539;
  wire signed [32-1:0] _reinterpretcast_src_540;
  assign _reinterpretcast_src_540 = _cond_data_481;
  wire signed [32-1:0] _reinterpretcast_data_540;
  assign _reinterpretcast_data_540 = _reinterpretcast_src_540;
  wire signed [32-1:0] _reinterpretcast_src_541;
  assign _reinterpretcast_src_541 = _cond_data_431;
  wire signed [32-1:0] _reinterpretcast_data_541;
  assign _reinterpretcast_data_541 = _reinterpretcast_src_541;
  wire signed [32-1:0] _reinterpretcast_src_542;
  assign _reinterpretcast_src_542 = _cond_data_461;
  wire signed [32-1:0] _reinterpretcast_data_542;
  assign _reinterpretcast_data_542 = _reinterpretcast_src_542;
  wire signed [32-1:0] _reinterpretcast_src_543;
  assign _reinterpretcast_src_543 = _cond_data_491;
  wire signed [32-1:0] _reinterpretcast_data_543;
  assign _reinterpretcast_data_543 = _reinterpretcast_src_543;
  wire signed [32-1:0] _reinterpretcast_src_544;
  assign _reinterpretcast_src_544 = _cond_data_441;
  wire signed [32-1:0] _reinterpretcast_data_544;
  assign _reinterpretcast_data_544 = _reinterpretcast_src_544;
  wire signed [32-1:0] _reinterpretcast_src_545;
  assign _reinterpretcast_src_545 = _cond_data_471;
  wire signed [32-1:0] _reinterpretcast_data_545;
  assign _reinterpretcast_data_545 = _reinterpretcast_src_545;
  wire signed [32-1:0] _reinterpretcast_src_546;
  assign _reinterpretcast_src_546 = _cond_data_501;
  wire signed [32-1:0] _reinterpretcast_data_546;
  assign _reinterpretcast_data_546 = _reinterpretcast_src_546;
  wire signed [32-1:0] _cond_data_620;
  assign _cond_data_620 = (__delay_data_875_pointer_601)? 1'sd0 : _reinterpretcast_data_538;
  wire signed [32-1:0] _cond_data_622;
  assign _cond_data_622 = (__delay_data_877_pointer_603)? 1'sd0 : _reinterpretcast_data_539;
  wire signed [32-1:0] _cond_data_624;
  assign _cond_data_624 = (__delay_data_879_pointer_605)? 1'sd0 : _reinterpretcast_data_540;
  wire signed [32-1:0] _cond_data_626;
  assign _cond_data_626 = (__delay_data_881_pointer_607)? 1'sd0 : _reinterpretcast_data_541;
  wire signed [32-1:0] _cond_data_628;
  assign _cond_data_628 = (__delay_data_883_pointer_609)? 1'sd0 : _reinterpretcast_data_542;
  wire signed [32-1:0] _cond_data_630;
  assign _cond_data_630 = (__delay_data_885_pointer_611)? 1'sd0 : _reinterpretcast_data_543;
  wire signed [32-1:0] _cond_data_632;
  assign _cond_data_632 = (__delay_data_887_pointer_613)? 1'sd0 : _reinterpretcast_data_544;
  wire signed [32-1:0] _cond_data_634;
  assign _cond_data_634 = (__delay_data_889_pointer_615)? 1'sd0 : _reinterpretcast_data_545;
  wire signed [32-1:0] _cond_data_636;
  assign _cond_data_636 = (__delay_data_891_pointer_617)? 1'sd0 : _reinterpretcast_data_546;
  reg signed [32-1:0] __variable_wdata_70;
  assign mul_3_x_data = __variable_wdata_70;
  reg signed [32-1:0] __variable_wdata_71;
  assign mul_3_y_data = __variable_wdata_71;
  reg [6-1:0] __variable_wdata_72;
  assign mul_3_rshift_data = __variable_wdata_72;
  assign _mul_3_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_3_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_3_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_91;
  assign mul_4_x_data = __variable_wdata_91;
  reg signed [32-1:0] __variable_wdata_92;
  assign mul_4_y_data = __variable_wdata_92;
  reg [6-1:0] __variable_wdata_93;
  assign mul_4_rshift_data = __variable_wdata_93;
  assign _mul_4_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_4_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_4_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_112;
  assign mul_5_x_data = __variable_wdata_112;
  reg signed [32-1:0] __variable_wdata_113;
  assign mul_5_y_data = __variable_wdata_113;
  reg [6-1:0] __variable_wdata_114;
  assign mul_5_rshift_data = __variable_wdata_114;
  assign _mul_5_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_5_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_5_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_133;
  assign mul_6_x_data = __variable_wdata_133;
  reg signed [32-1:0] __variable_wdata_134;
  assign mul_6_y_data = __variable_wdata_134;
  reg [6-1:0] __variable_wdata_135;
  assign mul_6_rshift_data = __variable_wdata_135;
  assign _mul_6_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_6_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_6_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_154;
  assign mul_7_x_data = __variable_wdata_154;
  reg signed [32-1:0] __variable_wdata_155;
  assign mul_7_y_data = __variable_wdata_155;
  reg [6-1:0] __variable_wdata_156;
  assign mul_7_rshift_data = __variable_wdata_156;
  assign _mul_7_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_7_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_7_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_175;
  assign mul_8_x_data = __variable_wdata_175;
  reg signed [32-1:0] __variable_wdata_176;
  assign mul_8_y_data = __variable_wdata_176;
  reg [6-1:0] __variable_wdata_177;
  assign mul_8_rshift_data = __variable_wdata_177;
  assign _mul_8_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_8_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_8_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_196;
  assign mul_9_x_data = __variable_wdata_196;
  reg signed [32-1:0] __variable_wdata_197;
  assign mul_9_y_data = __variable_wdata_197;
  reg [6-1:0] __variable_wdata_198;
  assign mul_9_rshift_data = __variable_wdata_198;
  assign _mul_9_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_9_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_9_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_217;
  assign mul_10_x_data = __variable_wdata_217;
  reg signed [32-1:0] __variable_wdata_218;
  assign mul_10_y_data = __variable_wdata_218;
  reg [6-1:0] __variable_wdata_219;
  assign mul_10_rshift_data = __variable_wdata_219;
  assign _mul_10_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_10_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_10_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_238;
  assign mul_11_x_data = __variable_wdata_238;
  reg signed [32-1:0] __variable_wdata_239;
  assign mul_11_y_data = __variable_wdata_239;
  reg [6-1:0] __variable_wdata_240;
  assign mul_11_rshift_data = __variable_wdata_240;
  assign _mul_11_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_11_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_11_stream_internal_oready;
  reg [1-1:0] __delay_data_894__delay_893__variable_264;
  reg [32-1:0] __delay_data_906_plus_822;
  reg [4-1:0] __delay_data_919__delay_918__variable_259;
  reg signed [32-1:0] __delay_data_932__delay_931_cond_280;
  reg signed [32-1:0] __delay_data_951__delay_950_cond_287;
  reg [32-1:0] __delay_data_970_plus_841;
  reg [1-1:0] __delay_data_895__delay_894__delay_893__variable_264;
  reg [32-1:0] __delay_data_907__delay_906_plus_822;
  reg [4-1:0] __delay_data_920__delay_919__delay_918__variable_259;
  reg signed [32-1:0] __delay_data_933__delay_932__delay_931_cond_280;
  reg signed [32-1:0] __delay_data_952__delay_951__delay_950_cond_287;
  reg [32-1:0] __delay_data_971__delay_970_plus_841;
  reg [1-1:0] __delay_data_896__delay_895__delay_894____variable_264;
  reg [32-1:0] __delay_data_908__delay_907__delay_906_plus_822;
  reg [4-1:0] __delay_data_921__delay_920__delay_919____variable_259;
  reg signed [32-1:0] __delay_data_934__delay_933__delay_932__delay_931_cond_280;
  reg signed [32-1:0] __delay_data_953__delay_952__delay_951__delay_950_cond_287;
  reg [32-1:0] __delay_data_972__delay_971__delay_970_plus_841;
  reg [1-1:0] __delay_data_897__delay_896__delay_895____variable_264;
  reg [32-1:0] __delay_data_909__delay_908__delay_907__delay_906_plus_822;
  reg [4-1:0] __delay_data_922__delay_921__delay_920____variable_259;
  reg signed [32-1:0] __delay_data_935__delay_934__delay_933__delay_932___cond_280;
  reg signed [32-1:0] __delay_data_954__delay_953__delay_952__delay_951___cond_287;
  reg [32-1:0] __delay_data_973__delay_972__delay_971__delay_970_plus_841;
  reg [1-1:0] __delay_data_898__delay_897__delay_896____variable_264;
  reg [32-1:0] __delay_data_910__delay_909__delay_908__delay_907___plus_822;
  reg [4-1:0] __delay_data_923__delay_922__delay_921____variable_259;
  reg signed [32-1:0] __delay_data_936__delay_935__delay_934__delay_933___cond_280;
  reg signed [32-1:0] __delay_data_955__delay_954__delay_953__delay_952___cond_287;
  reg [32-1:0] __delay_data_974__delay_973__delay_972__delay_971___plus_841;
  reg [1-1:0] __delay_data_899__delay_898__delay_897____variable_264;
  reg [32-1:0] __delay_data_911__delay_910__delay_909__delay_908___plus_822;
  reg [4-1:0] __delay_data_924__delay_923__delay_922____variable_259;
  reg signed [32-1:0] __delay_data_937__delay_936__delay_935__delay_934___cond_280;
  reg signed [32-1:0] __delay_data_956__delay_955__delay_954__delay_953___cond_287;
  reg [32-1:0] __delay_data_975__delay_974__delay_973__delay_972___plus_841;
  reg [1-1:0] __delay_data_900__delay_899__delay_898____variable_264;
  reg [32-1:0] __delay_data_912__delay_911__delay_910__delay_909___plus_822;
  reg [4-1:0] __delay_data_925__delay_924__delay_923____variable_259;
  reg signed [32-1:0] __delay_data_938__delay_937__delay_936__delay_935___cond_280;
  reg signed [32-1:0] __delay_data_957__delay_956__delay_955__delay_954___cond_287;
  reg [32-1:0] __delay_data_976__delay_975__delay_974__delay_973___plus_841;
  reg [1-1:0] __delay_data_901__delay_900__delay_899____variable_264;
  reg [32-1:0] __delay_data_913__delay_912__delay_911__delay_910___plus_822;
  reg [4-1:0] __delay_data_926__delay_925__delay_924____variable_259;
  reg signed [32-1:0] __delay_data_939__delay_938__delay_937__delay_936___cond_280;
  reg signed [32-1:0] __delay_data_958__delay_957__delay_956__delay_955___cond_287;
  reg [32-1:0] __delay_data_977__delay_976__delay_975__delay_974___plus_841;
  reg [1-1:0] __delay_data_902__delay_901__delay_900____variable_264;
  reg [32-1:0] __delay_data_914__delay_913__delay_912__delay_911___plus_822;
  reg [4-1:0] __delay_data_927__delay_926__delay_925____variable_259;
  reg signed [32-1:0] __delay_data_940__delay_939__delay_938__delay_937___cond_280;
  reg signed [32-1:0] __delay_data_959__delay_958__delay_957__delay_956___cond_287;
  reg [32-1:0] __delay_data_978__delay_977__delay_976__delay_975___plus_841;
  wire signed [32-1:0] __substreamoutput_data_655;
  assign __substreamoutput_data_655 = mul_3_z_data;
  wire signed [32-1:0] __substreamoutput_data_674;
  assign __substreamoutput_data_674 = mul_4_z_data;
  wire signed [32-1:0] __substreamoutput_data_693;
  assign __substreamoutput_data_693 = mul_5_z_data;
  wire signed [32-1:0] __substreamoutput_data_712;
  assign __substreamoutput_data_712 = mul_6_z_data;
  wire signed [32-1:0] __substreamoutput_data_731;
  assign __substreamoutput_data_731 = mul_7_z_data;
  wire signed [32-1:0] __substreamoutput_data_750;
  assign __substreamoutput_data_750 = mul_8_z_data;
  wire signed [32-1:0] __substreamoutput_data_769;
  assign __substreamoutput_data_769 = mul_9_z_data;
  wire signed [32-1:0] __substreamoutput_data_788;
  assign __substreamoutput_data_788 = mul_10_z_data;
  wire signed [32-1:0] __substreamoutput_data_807;
  assign __substreamoutput_data_807 = mul_11_z_data;
  reg signed [32-1:0] __variable_wdata_22;
  assign add_tree_1_var0_data = __variable_wdata_22;
  reg signed [32-1:0] __variable_wdata_23;
  assign add_tree_1_var1_data = __variable_wdata_23;
  reg signed [32-1:0] __variable_wdata_24;
  assign add_tree_1_var2_data = __variable_wdata_24;
  reg signed [32-1:0] __variable_wdata_25;
  assign add_tree_1_var3_data = __variable_wdata_25;
  reg signed [32-1:0] __variable_wdata_26;
  assign add_tree_1_var4_data = __variable_wdata_26;
  reg signed [32-1:0] __variable_wdata_27;
  assign add_tree_1_var5_data = __variable_wdata_27;
  reg signed [32-1:0] __variable_wdata_28;
  assign add_tree_1_var6_data = __variable_wdata_28;
  reg signed [32-1:0] __variable_wdata_29;
  assign add_tree_1_var7_data = __variable_wdata_29;
  reg signed [32-1:0] __variable_wdata_30;
  assign add_tree_1_var8_data = __variable_wdata_30;
  assign _add_tree_1_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _add_tree_1_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _add_tree_1_stream_internal_oready;
  reg [1-1:0] __delay_data_903__delay_902__delay_901____variable_264;
  reg [32-1:0] __delay_data_915__delay_914__delay_913__delay_912___plus_822;
  reg [4-1:0] __delay_data_928__delay_927__delay_926____variable_259;
  reg signed [32-1:0] __delay_data_941__delay_940__delay_939__delay_938___cond_280;
  reg signed [32-1:0] __delay_data_960__delay_959__delay_958__delay_957___cond_287;
  reg [32-1:0] __delay_data_979__delay_978__delay_977__delay_976___plus_841;
  reg [1-1:0] __delay_data_904__delay_903__delay_902____variable_264;
  reg [32-1:0] __delay_data_916__delay_915__delay_914__delay_913___plus_822;
  reg [4-1:0] __delay_data_929__delay_928__delay_927____variable_259;
  reg signed [32-1:0] __delay_data_942__delay_941__delay_940__delay_939___cond_280;
  reg signed [32-1:0] __delay_data_961__delay_960__delay_959__delay_958___cond_287;
  reg [32-1:0] __delay_data_980__delay_979__delay_978__delay_977___plus_841;
  reg [1-1:0] __delay_data_905__delay_904__delay_903____variable_264;
  reg [32-1:0] __delay_data_917__delay_916__delay_915__delay_914___plus_822;
  reg [4-1:0] __delay_data_930__delay_929__delay_928____variable_259;
  reg signed [32-1:0] __delay_data_943__delay_942__delay_941__delay_940___cond_280;
  reg signed [32-1:0] __delay_data_962__delay_961__delay_960__delay_959___cond_287;
  reg [32-1:0] __delay_data_981__delay_980__delay_979__delay_978___plus_841;
  wire signed [32-1:0] __substreamoutput_data_809;
  assign __substreamoutput_data_809 = add_tree_1_sum_data;
  reg [1-1:0] __variable_wdata_15;
  assign acc_0__reduce_reset_data = __variable_wdata_15;
  reg signed [32-1:0] __variable_wdata_0;
  assign acc_0_x_data = __variable_wdata_0;
  reg [6-1:0] __variable_wdata_1;
  assign acc_0_rshift_data = __variable_wdata_1;
  reg [32-1:0] __variable_wdata_2;
  assign acc_0_size_data = __variable_wdata_2;
  assign _acc_0_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _acc_0_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _acc_0_stream_internal_oready;
  reg signed [32-1:0] __delay_data_944__delay_943__delay_942__delay_941___cond_280;
  reg signed [32-1:0] __delay_data_963__delay_962__delay_961__delay_960___cond_287;
  reg [32-1:0] __delay_data_982__delay_981__delay_980__delay_979___plus_841;
  reg signed [32-1:0] __delay_data_945__delay_944__delay_943__delay_942___cond_280;
  reg signed [32-1:0] __delay_data_964__delay_963__delay_962__delay_961___cond_287;
  reg [32-1:0] __delay_data_983__delay_982__delay_981__delay_980___plus_841;
  reg signed [32-1:0] __delay_data_946__delay_945__delay_944__delay_943___cond_280;
  reg signed [32-1:0] __delay_data_965__delay_964__delay_963__delay_962___cond_287;
  reg [32-1:0] __delay_data_984__delay_983__delay_982__delay_981___plus_841;
  reg signed [32-1:0] __delay_data_947__delay_946__delay_945__delay_944___cond_280;
  reg signed [32-1:0] __delay_data_966__delay_965__delay_964__delay_963___cond_287;
  reg [32-1:0] __delay_data_985__delay_984__delay_983__delay_982___plus_841;
  reg signed [32-1:0] __delay_data_948__delay_947__delay_946__delay_945___cond_280;
  reg signed [32-1:0] __delay_data_967__delay_966__delay_965__delay_964___cond_287;
  reg [32-1:0] __delay_data_986__delay_985__delay_984__delay_983___plus_841;
  reg signed [32-1:0] __delay_data_949__delay_948__delay_947__delay_946___cond_280;
  reg signed [32-1:0] __delay_data_968__delay_967__delay_966__delay_965___cond_287;
  reg [32-1:0] __delay_data_987__delay_986__delay_985__delay_984___plus_841;
  wire signed [32-1:0] __substreamoutput_data_823;
  assign __substreamoutput_data_823 = acc_0_sum_data;
  wire [1-1:0] __substreamoutput_data_824;
  assign __substreamoutput_data_824 = acc_0_valid_data;
  reg signed [32-1:0] _plus_data_825;
  reg signed [32-1:0] __delay_data_969__delay_968__delay_967__delay_966___cond_287;
  reg [32-1:0] __delay_data_988__delay_987__delay_986__delay_985___plus_841;
  reg [1-1:0] __delay_data_989__substreamoutput_824;
  reg signed [32-1:0] __variable_wdata_36;
  assign mul_rshift_round_clip_2_x_data = __variable_wdata_36;
  reg signed [32-1:0] __variable_wdata_37;
  assign mul_rshift_round_clip_2_y_data = __variable_wdata_37;
  reg [6-1:0] __variable_wdata_38;
  assign mul_rshift_round_clip_2_rshift_data = __variable_wdata_38;
  assign _mul_rshift_round_clip_2_is_root = ((_stream_conv2d_2_busy)? 0 : 1) && 1;
  assign _mul_rshift_round_clip_2_stream_oready = ((_stream_conv2d_2_busy)? _stream_conv2d_2_stream_oready : 1) && _mul_rshift_round_clip_2_stream_internal_oready;
  assign _stream_conv2d_2_stream_internal_oready = ((_stream_conv2d_2_busy)? _mul_rshift_round_clip_2_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _acc_0_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _add_tree_1_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_11_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_10_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_9_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_8_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_7_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_6_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_5_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_4_stream_internal_oready : 1) && (((_stream_conv2d_2_busy)? _mul_3_stream_internal_oready : 1) && 1)))))))))));
  reg [1-1:0] __delay_data_990__delay_989__substreamoutput_824;
  reg [1-1:0] __delay_data_991__delay_990__delay_989__substreamoutput_824;
  reg [1-1:0] __delay_data_992__delay_991__delay_990____substreamoutput_824;
  reg [1-1:0] __delay_data_993__delay_992__delay_991____substreamoutput_824;
  reg [1-1:0] __delay_data_994__delay_993__delay_992____substreamoutput_824;
  reg [1-1:0] __delay_data_995__delay_994__delay_993____substreamoutput_824;
  reg [1-1:0] __delay_data_996__delay_995__delay_994____substreamoutput_824;
  reg [1-1:0] __delay_data_997__delay_996__delay_995____substreamoutput_824;
  reg [1-1:0] __delay_data_998__delay_997__delay_996____substreamoutput_824;
  wire signed [32-1:0] __substreamoutput_data_842;
  assign __substreamoutput_data_842 = mul_rshift_round_clip_2_z_data;
  wire signed [32-1:0] _reinterpretcast_src_843;
  assign _reinterpretcast_src_843 = __substreamoutput_data_842;
  wire signed [32-1:0] _reinterpretcast_data_843;
  assign _reinterpretcast_data_843 = _reinterpretcast_src_843;
  wire signed [32-1:0] stream_conv2d_2_sink_50_data;
  assign stream_conv2d_2_sink_50_data = _reinterpretcast_data_843;
  wire [1-1:0] stream_conv2d_2_sink_51_data;
  assign stream_conv2d_2_sink_51_data = __delay_data_998__delay_997__delay_996____substreamoutput_824;
  wire _set_flag_177;
  assign _set_flag_177 = conv2d_2_comp_fsm == 3;
  reg [4-1:0] __variable_wdata_259;
  assign stream_conv2d_2_parameter_0_data = __variable_wdata_259;
  wire _set_flag_178;
  assign _set_flag_178 = conv2d_2_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_260;
  assign stream_conv2d_2_parameter_1_data = __variable_wdata_260;
  wire _set_flag_179;
  assign _set_flag_179 = conv2d_2_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_261;
  assign stream_conv2d_2_parameter_2_data = __variable_wdata_261;
  wire _set_flag_180;
  assign _set_flag_180 = conv2d_2_comp_fsm == 3;
  reg [9-1:0] __variable_wdata_262;
  assign stream_conv2d_2_parameter_3_data = __variable_wdata_262;
  wire _set_flag_181;
  assign _set_flag_181 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_263;
  assign stream_conv2d_2_parameter_4_data = __variable_wdata_263;
  wire _set_flag_182;
  assign _set_flag_182 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_274;
  assign stream_conv2d_2_parameter_6_data = __variable_wdata_274;
  wire _set_flag_183;
  assign _set_flag_183 = conv2d_2_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_275;
  assign stream_conv2d_2_source_7_data = __variable_wdata_275;
  wire _set_flag_184;
  assign _set_flag_184 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_281;
  assign stream_conv2d_2_parameter_8_data = __variable_wdata_281;
  wire _set_flag_185;
  assign _set_flag_185 = conv2d_2_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_282;
  assign stream_conv2d_2_source_9_data = __variable_wdata_282;
  wire _set_flag_186;
  assign _set_flag_186 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_288;
  assign stream_conv2d_2_parameter_10_data = __variable_wdata_288;
  wire _set_flag_187;
  assign _set_flag_187 = conv2d_2_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_289;
  assign stream_conv2d_2_source_11_data = __variable_wdata_289;
  wire _set_flag_188;
  assign _set_flag_188 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_295;
  assign stream_conv2d_2_parameter_12_data = __variable_wdata_295;
  wire _set_flag_189;
  assign _set_flag_189 = conv2d_2_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_296;
  assign stream_conv2d_2_source_13_data = __variable_wdata_296;
  wire _set_flag_190;
  assign _set_flag_190 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_302;
  assign stream_conv2d_2_parameter_14_data = __variable_wdata_302;
  wire _set_flag_191;
  assign _set_flag_191 = conv2d_2_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_303;
  assign stream_conv2d_2_source_15_data = __variable_wdata_303;
  wire _set_flag_192;
  assign _set_flag_192 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_309;
  assign stream_conv2d_2_parameter_16_data = __variable_wdata_309;
  wire _set_flag_193;
  assign _set_flag_193 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_310;
  assign stream_conv2d_2_parameter_17_data = __variable_wdata_310;
  wire _set_flag_194;
  assign _set_flag_194 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_311;
  assign stream_conv2d_2_parameter_18_data = __variable_wdata_311;
  wire _set_flag_195;
  assign _set_flag_195 = conv2d_2_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_312;
  assign stream_conv2d_2_parameter_19_data = __variable_wdata_312;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_20_pat_stride_buf_3;
  wire _set_flag_196;
  assign _set_flag_196 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id10_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_20_source_ram_renable && (_stream_conv2d_2_source_20_source_sel == 1))? _stream_conv2d_2_source_20_source_ram_raddr : 'hx;
  assign ram_w32_l128_id10_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_20_source_ram_renable && (_stream_conv2d_2_source_20_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_197 = 1;
  wire [_tmp_197-1:0] _tmp_198;
  assign _tmp_198 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_20_source_ram_renable && (_stream_conv2d_2_source_20_source_sel == 1);
  reg [_tmp_197-1:0] __tmp_198_1;
  assign _stream_conv2d_2_source_20_source_ram_rdata = (_stream_conv2d_2_source_20_source_sel == 1)? ram_w32_l128_id10_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_313;
  assign stream_conv2d_2_source_20_data = __variable_wdata_313;
  reg [32-1:0] _stream_conv2d_2_source_20_source_pat_fsm_0;
  localparam _stream_conv2d_2_source_20_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_20_source_pat_all_offset;
  assign _stream_conv2d_2_source_20_source_pat_all_offset = _stream_conv2d_2_source_20_source_offset_buf + _source_stream_conv2d_2_source_20_pat_cur_offset_0 + _source_stream_conv2d_2_source_20_pat_cur_offset_1 + _source_stream_conv2d_2_source_20_pat_cur_offset_2 + _source_stream_conv2d_2_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_21_pat_stride_buf_3;
  wire _set_flag_199;
  assign _set_flag_199 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id11_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_21_source_ram_renable && (_stream_conv2d_2_source_21_source_sel == 2))? _stream_conv2d_2_source_21_source_ram_raddr : 'hx;
  assign ram_w32_l128_id11_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_21_source_ram_renable && (_stream_conv2d_2_source_21_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_200 = 1;
  wire [_tmp_200-1:0] _tmp_201;
  assign _tmp_201 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_21_source_ram_renable && (_stream_conv2d_2_source_21_source_sel == 2);
  reg [_tmp_200-1:0] __tmp_201_1;
  assign _stream_conv2d_2_source_21_source_ram_rdata = (_stream_conv2d_2_source_21_source_sel == 2)? ram_w32_l128_id11_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_314;
  assign stream_conv2d_2_source_21_data = __variable_wdata_314;
  reg [32-1:0] _stream_conv2d_2_source_21_source_pat_fsm_1;
  localparam _stream_conv2d_2_source_21_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_21_source_pat_all_offset;
  assign _stream_conv2d_2_source_21_source_pat_all_offset = _stream_conv2d_2_source_21_source_offset_buf + _source_stream_conv2d_2_source_21_pat_cur_offset_0 + _source_stream_conv2d_2_source_21_pat_cur_offset_1 + _source_stream_conv2d_2_source_21_pat_cur_offset_2 + _source_stream_conv2d_2_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_22_pat_stride_buf_3;
  wire _set_flag_202;
  assign _set_flag_202 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id12_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_22_source_ram_renable && (_stream_conv2d_2_source_22_source_sel == 3))? _stream_conv2d_2_source_22_source_ram_raddr : 'hx;
  assign ram_w32_l128_id12_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_22_source_ram_renable && (_stream_conv2d_2_source_22_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_203 = 1;
  wire [_tmp_203-1:0] _tmp_204;
  assign _tmp_204 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_22_source_ram_renable && (_stream_conv2d_2_source_22_source_sel == 3);
  reg [_tmp_203-1:0] __tmp_204_1;
  assign _stream_conv2d_2_source_22_source_ram_rdata = (_stream_conv2d_2_source_22_source_sel == 3)? ram_w32_l128_id12_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_315;
  assign stream_conv2d_2_source_22_data = __variable_wdata_315;
  reg [32-1:0] _stream_conv2d_2_source_22_source_pat_fsm_2;
  localparam _stream_conv2d_2_source_22_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_22_source_pat_all_offset;
  assign _stream_conv2d_2_source_22_source_pat_all_offset = _stream_conv2d_2_source_22_source_offset_buf + _source_stream_conv2d_2_source_22_pat_cur_offset_0 + _source_stream_conv2d_2_source_22_pat_cur_offset_1 + _source_stream_conv2d_2_source_22_pat_cur_offset_2 + _source_stream_conv2d_2_source_22_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_23_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_23_pat_stride_buf_3;
  wire _set_flag_205;
  assign _set_flag_205 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id13_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_23_source_ram_renable && (_stream_conv2d_2_source_23_source_sel == 4))? _stream_conv2d_2_source_23_source_ram_raddr : 'hx;
  assign ram_w32_l128_id13_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_23_source_ram_renable && (_stream_conv2d_2_source_23_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_206 = 1;
  wire [_tmp_206-1:0] _tmp_207;
  assign _tmp_207 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_23_source_ram_renable && (_stream_conv2d_2_source_23_source_sel == 4);
  reg [_tmp_206-1:0] __tmp_207_1;
  assign _stream_conv2d_2_source_23_source_ram_rdata = (_stream_conv2d_2_source_23_source_sel == 4)? ram_w32_l128_id13_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_316;
  assign stream_conv2d_2_source_23_data = __variable_wdata_316;
  reg [32-1:0] _stream_conv2d_2_source_23_source_pat_fsm_3;
  localparam _stream_conv2d_2_source_23_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_23_source_pat_all_offset;
  assign _stream_conv2d_2_source_23_source_pat_all_offset = _stream_conv2d_2_source_23_source_offset_buf + _source_stream_conv2d_2_source_23_pat_cur_offset_0 + _source_stream_conv2d_2_source_23_pat_cur_offset_1 + _source_stream_conv2d_2_source_23_pat_cur_offset_2 + _source_stream_conv2d_2_source_23_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_24_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_24_pat_stride_buf_3;
  wire _set_flag_208;
  assign _set_flag_208 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id14_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_24_source_ram_renable && (_stream_conv2d_2_source_24_source_sel == 5))? _stream_conv2d_2_source_24_source_ram_raddr : 'hx;
  assign ram_w32_l128_id14_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_24_source_ram_renable && (_stream_conv2d_2_source_24_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_209 = 1;
  wire [_tmp_209-1:0] _tmp_210;
  assign _tmp_210 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_24_source_ram_renable && (_stream_conv2d_2_source_24_source_sel == 5);
  reg [_tmp_209-1:0] __tmp_210_1;
  assign _stream_conv2d_2_source_24_source_ram_rdata = (_stream_conv2d_2_source_24_source_sel == 5)? ram_w32_l128_id14_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_317;
  assign stream_conv2d_2_source_24_data = __variable_wdata_317;
  reg [32-1:0] _stream_conv2d_2_source_24_source_pat_fsm_4;
  localparam _stream_conv2d_2_source_24_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_24_source_pat_all_offset;
  assign _stream_conv2d_2_source_24_source_pat_all_offset = _stream_conv2d_2_source_24_source_offset_buf + _source_stream_conv2d_2_source_24_pat_cur_offset_0 + _source_stream_conv2d_2_source_24_pat_cur_offset_1 + _source_stream_conv2d_2_source_24_pat_cur_offset_2 + _source_stream_conv2d_2_source_24_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_25_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_25_pat_stride_buf_3;
  wire _set_flag_211;
  assign _set_flag_211 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id15_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_25_source_ram_renable && (_stream_conv2d_2_source_25_source_sel == 6))? _stream_conv2d_2_source_25_source_ram_raddr : 'hx;
  assign ram_w32_l128_id15_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_25_source_ram_renable && (_stream_conv2d_2_source_25_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_212 = 1;
  wire [_tmp_212-1:0] _tmp_213;
  assign _tmp_213 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_25_source_ram_renable && (_stream_conv2d_2_source_25_source_sel == 6);
  reg [_tmp_212-1:0] __tmp_213_1;
  assign _stream_conv2d_2_source_25_source_ram_rdata = (_stream_conv2d_2_source_25_source_sel == 6)? ram_w32_l128_id15_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_318;
  assign stream_conv2d_2_source_25_data = __variable_wdata_318;
  reg [32-1:0] _stream_conv2d_2_source_25_source_pat_fsm_5;
  localparam _stream_conv2d_2_source_25_source_pat_fsm_5_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_25_source_pat_all_offset;
  assign _stream_conv2d_2_source_25_source_pat_all_offset = _stream_conv2d_2_source_25_source_offset_buf + _source_stream_conv2d_2_source_25_pat_cur_offset_0 + _source_stream_conv2d_2_source_25_pat_cur_offset_1 + _source_stream_conv2d_2_source_25_pat_cur_offset_2 + _source_stream_conv2d_2_source_25_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_26_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_26_pat_stride_buf_3;
  wire _set_flag_214;
  assign _set_flag_214 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id16_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_26_source_ram_renable && (_stream_conv2d_2_source_26_source_sel == 7))? _stream_conv2d_2_source_26_source_ram_raddr : 'hx;
  assign ram_w32_l128_id16_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_26_source_ram_renable && (_stream_conv2d_2_source_26_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_215 = 1;
  wire [_tmp_215-1:0] _tmp_216;
  assign _tmp_216 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_26_source_ram_renable && (_stream_conv2d_2_source_26_source_sel == 7);
  reg [_tmp_215-1:0] __tmp_216_1;
  assign _stream_conv2d_2_source_26_source_ram_rdata = (_stream_conv2d_2_source_26_source_sel == 7)? ram_w32_l128_id16_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_319;
  assign stream_conv2d_2_source_26_data = __variable_wdata_319;
  reg [32-1:0] _stream_conv2d_2_source_26_source_pat_fsm_6;
  localparam _stream_conv2d_2_source_26_source_pat_fsm_6_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_26_source_pat_all_offset;
  assign _stream_conv2d_2_source_26_source_pat_all_offset = _stream_conv2d_2_source_26_source_offset_buf + _source_stream_conv2d_2_source_26_pat_cur_offset_0 + _source_stream_conv2d_2_source_26_pat_cur_offset_1 + _source_stream_conv2d_2_source_26_pat_cur_offset_2 + _source_stream_conv2d_2_source_26_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_27_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_27_pat_stride_buf_3;
  wire _set_flag_217;
  assign _set_flag_217 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id17_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_27_source_ram_renable && (_stream_conv2d_2_source_27_source_sel == 8))? _stream_conv2d_2_source_27_source_ram_raddr : 'hx;
  assign ram_w32_l128_id17_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_27_source_ram_renable && (_stream_conv2d_2_source_27_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_218 = 1;
  wire [_tmp_218-1:0] _tmp_219;
  assign _tmp_219 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_27_source_ram_renable && (_stream_conv2d_2_source_27_source_sel == 8);
  reg [_tmp_218-1:0] __tmp_219_1;
  assign _stream_conv2d_2_source_27_source_ram_rdata = (_stream_conv2d_2_source_27_source_sel == 8)? ram_w32_l128_id17_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_320;
  assign stream_conv2d_2_source_27_data = __variable_wdata_320;
  reg [32-1:0] _stream_conv2d_2_source_27_source_pat_fsm_7;
  localparam _stream_conv2d_2_source_27_source_pat_fsm_7_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_27_source_pat_all_offset;
  assign _stream_conv2d_2_source_27_source_pat_all_offset = _stream_conv2d_2_source_27_source_offset_buf + _source_stream_conv2d_2_source_27_pat_cur_offset_0 + _source_stream_conv2d_2_source_27_pat_cur_offset_1 + _source_stream_conv2d_2_source_27_pat_cur_offset_2 + _source_stream_conv2d_2_source_27_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_28_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_28_pat_stride_buf_3;
  wire _set_flag_220;
  assign _set_flag_220 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id18_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_28_source_ram_renable && (_stream_conv2d_2_source_28_source_sel == 9))? _stream_conv2d_2_source_28_source_ram_raddr : 'hx;
  assign ram_w32_l128_id18_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_28_source_ram_renable && (_stream_conv2d_2_source_28_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_221 = 1;
  wire [_tmp_221-1:0] _tmp_222;
  assign _tmp_222 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_28_source_ram_renable && (_stream_conv2d_2_source_28_source_sel == 9);
  reg [_tmp_221-1:0] __tmp_222_1;
  assign _stream_conv2d_2_source_28_source_ram_rdata = (_stream_conv2d_2_source_28_source_sel == 9)? ram_w32_l128_id18_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_321;
  assign stream_conv2d_2_source_28_data = __variable_wdata_321;
  reg [32-1:0] _stream_conv2d_2_source_28_source_pat_fsm_8;
  localparam _stream_conv2d_2_source_28_source_pat_fsm_8_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_28_source_pat_all_offset;
  assign _stream_conv2d_2_source_28_source_pat_all_offset = _stream_conv2d_2_source_28_source_offset_buf + _source_stream_conv2d_2_source_28_pat_cur_offset_0 + _source_stream_conv2d_2_source_28_pat_cur_offset_1 + _source_stream_conv2d_2_source_28_pat_cur_offset_2 + _source_stream_conv2d_2_source_28_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_29_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_29_pat_stride_buf_3;
  wire _set_flag_223;
  assign _set_flag_223 = conv2d_2_comp_fsm == 3;
  localparam _tmp_224 = 1;
  wire [_tmp_224-1:0] _tmp_225;
  assign _tmp_225 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_29_source_ram_renable && (_stream_conv2d_2_source_29_source_sel == 10);
  reg [_tmp_224-1:0] __tmp_225_1;
  assign _stream_conv2d_2_source_29_source_ram_rdata = (_stream_conv2d_2_source_29_source_sel == 10)? ram_w32_l128_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_547;
  assign stream_conv2d_2_source_29_data = __variable_wdata_547;
  reg [32-1:0] _stream_conv2d_2_source_29_source_pat_fsm_9;
  localparam _stream_conv2d_2_source_29_source_pat_fsm_9_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_29_source_pat_all_offset;
  assign _stream_conv2d_2_source_29_source_pat_all_offset = _stream_conv2d_2_source_29_source_offset_buf + _source_stream_conv2d_2_source_29_pat_cur_offset_0 + _source_stream_conv2d_2_source_29_pat_cur_offset_1 + _source_stream_conv2d_2_source_29_pat_cur_offset_2 + _source_stream_conv2d_2_source_29_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_30_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_30_pat_stride_buf_3;
  wire _set_flag_226;
  assign _set_flag_226 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id2_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_30_source_ram_renable && (_stream_conv2d_2_source_30_source_sel == 11))? _stream_conv2d_2_source_30_source_ram_raddr : 'hx;
  assign ram_w32_l128_id2_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_30_source_ram_renable && (_stream_conv2d_2_source_30_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_227 = 1;
  wire [_tmp_227-1:0] _tmp_228;
  assign _tmp_228 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_30_source_ram_renable && (_stream_conv2d_2_source_30_source_sel == 11);
  reg [_tmp_227-1:0] __tmp_228_1;
  assign _stream_conv2d_2_source_30_source_ram_rdata = (_stream_conv2d_2_source_30_source_sel == 11)? ram_w32_l128_id2_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_548;
  assign stream_conv2d_2_source_30_data = __variable_wdata_548;
  reg [32-1:0] _stream_conv2d_2_source_30_source_pat_fsm_10;
  localparam _stream_conv2d_2_source_30_source_pat_fsm_10_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_30_source_pat_all_offset;
  assign _stream_conv2d_2_source_30_source_pat_all_offset = _stream_conv2d_2_source_30_source_offset_buf + _source_stream_conv2d_2_source_30_pat_cur_offset_0 + _source_stream_conv2d_2_source_30_pat_cur_offset_1 + _source_stream_conv2d_2_source_30_pat_cur_offset_2 + _source_stream_conv2d_2_source_30_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_31_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_31_pat_stride_buf_3;
  wire _set_flag_229;
  assign _set_flag_229 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id3_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_31_source_ram_renable && (_stream_conv2d_2_source_31_source_sel == 12))? _stream_conv2d_2_source_31_source_ram_raddr : 'hx;
  assign ram_w32_l128_id3_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_31_source_ram_renable && (_stream_conv2d_2_source_31_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_230 = 1;
  wire [_tmp_230-1:0] _tmp_231;
  assign _tmp_231 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_31_source_ram_renable && (_stream_conv2d_2_source_31_source_sel == 12);
  reg [_tmp_230-1:0] __tmp_231_1;
  assign _stream_conv2d_2_source_31_source_ram_rdata = (_stream_conv2d_2_source_31_source_sel == 12)? ram_w32_l128_id3_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_549;
  assign stream_conv2d_2_source_31_data = __variable_wdata_549;
  reg [32-1:0] _stream_conv2d_2_source_31_source_pat_fsm_11;
  localparam _stream_conv2d_2_source_31_source_pat_fsm_11_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_31_source_pat_all_offset;
  assign _stream_conv2d_2_source_31_source_pat_all_offset = _stream_conv2d_2_source_31_source_offset_buf + _source_stream_conv2d_2_source_31_pat_cur_offset_0 + _source_stream_conv2d_2_source_31_pat_cur_offset_1 + _source_stream_conv2d_2_source_31_pat_cur_offset_2 + _source_stream_conv2d_2_source_31_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_32_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_32_pat_stride_buf_3;
  wire _set_flag_232;
  assign _set_flag_232 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id4_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_32_source_ram_renable && (_stream_conv2d_2_source_32_source_sel == 13))? _stream_conv2d_2_source_32_source_ram_raddr : 'hx;
  assign ram_w32_l128_id4_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_32_source_ram_renable && (_stream_conv2d_2_source_32_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_233 = 1;
  wire [_tmp_233-1:0] _tmp_234;
  assign _tmp_234 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_32_source_ram_renable && (_stream_conv2d_2_source_32_source_sel == 13);
  reg [_tmp_233-1:0] __tmp_234_1;
  assign _stream_conv2d_2_source_32_source_ram_rdata = (_stream_conv2d_2_source_32_source_sel == 13)? ram_w32_l128_id4_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_550;
  assign stream_conv2d_2_source_32_data = __variable_wdata_550;
  reg [32-1:0] _stream_conv2d_2_source_32_source_pat_fsm_12;
  localparam _stream_conv2d_2_source_32_source_pat_fsm_12_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_32_source_pat_all_offset;
  assign _stream_conv2d_2_source_32_source_pat_all_offset = _stream_conv2d_2_source_32_source_offset_buf + _source_stream_conv2d_2_source_32_pat_cur_offset_0 + _source_stream_conv2d_2_source_32_pat_cur_offset_1 + _source_stream_conv2d_2_source_32_pat_cur_offset_2 + _source_stream_conv2d_2_source_32_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_33_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_33_pat_stride_buf_3;
  wire _set_flag_235;
  assign _set_flag_235 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id5_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_33_source_ram_renable && (_stream_conv2d_2_source_33_source_sel == 14))? _stream_conv2d_2_source_33_source_ram_raddr : 'hx;
  assign ram_w32_l128_id5_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_33_source_ram_renable && (_stream_conv2d_2_source_33_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_236 = 1;
  wire [_tmp_236-1:0] _tmp_237;
  assign _tmp_237 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_33_source_ram_renable && (_stream_conv2d_2_source_33_source_sel == 14);
  reg [_tmp_236-1:0] __tmp_237_1;
  assign _stream_conv2d_2_source_33_source_ram_rdata = (_stream_conv2d_2_source_33_source_sel == 14)? ram_w32_l128_id5_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_551;
  assign stream_conv2d_2_source_33_data = __variable_wdata_551;
  reg [32-1:0] _stream_conv2d_2_source_33_source_pat_fsm_13;
  localparam _stream_conv2d_2_source_33_source_pat_fsm_13_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_33_source_pat_all_offset;
  assign _stream_conv2d_2_source_33_source_pat_all_offset = _stream_conv2d_2_source_33_source_offset_buf + _source_stream_conv2d_2_source_33_pat_cur_offset_0 + _source_stream_conv2d_2_source_33_pat_cur_offset_1 + _source_stream_conv2d_2_source_33_pat_cur_offset_2 + _source_stream_conv2d_2_source_33_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_34_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_34_pat_stride_buf_3;
  wire _set_flag_238;
  assign _set_flag_238 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id6_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_34_source_ram_renable && (_stream_conv2d_2_source_34_source_sel == 15))? _stream_conv2d_2_source_34_source_ram_raddr : 'hx;
  assign ram_w32_l128_id6_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_34_source_ram_renable && (_stream_conv2d_2_source_34_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_239 = 1;
  wire [_tmp_239-1:0] _tmp_240;
  assign _tmp_240 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_34_source_ram_renable && (_stream_conv2d_2_source_34_source_sel == 15);
  reg [_tmp_239-1:0] __tmp_240_1;
  assign _stream_conv2d_2_source_34_source_ram_rdata = (_stream_conv2d_2_source_34_source_sel == 15)? ram_w32_l128_id6_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_552;
  assign stream_conv2d_2_source_34_data = __variable_wdata_552;
  reg [32-1:0] _stream_conv2d_2_source_34_source_pat_fsm_14;
  localparam _stream_conv2d_2_source_34_source_pat_fsm_14_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_34_source_pat_all_offset;
  assign _stream_conv2d_2_source_34_source_pat_all_offset = _stream_conv2d_2_source_34_source_offset_buf + _source_stream_conv2d_2_source_34_pat_cur_offset_0 + _source_stream_conv2d_2_source_34_pat_cur_offset_1 + _source_stream_conv2d_2_source_34_pat_cur_offset_2 + _source_stream_conv2d_2_source_34_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_35_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_35_pat_stride_buf_3;
  wire _set_flag_241;
  assign _set_flag_241 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id7_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_35_source_ram_renable && (_stream_conv2d_2_source_35_source_sel == 16))? _stream_conv2d_2_source_35_source_ram_raddr : 'hx;
  assign ram_w32_l128_id7_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_35_source_ram_renable && (_stream_conv2d_2_source_35_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_242 = 1;
  wire [_tmp_242-1:0] _tmp_243;
  assign _tmp_243 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_35_source_ram_renable && (_stream_conv2d_2_source_35_source_sel == 16);
  reg [_tmp_242-1:0] __tmp_243_1;
  assign _stream_conv2d_2_source_35_source_ram_rdata = (_stream_conv2d_2_source_35_source_sel == 16)? ram_w32_l128_id7_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_553;
  assign stream_conv2d_2_source_35_data = __variable_wdata_553;
  reg [32-1:0] _stream_conv2d_2_source_35_source_pat_fsm_15;
  localparam _stream_conv2d_2_source_35_source_pat_fsm_15_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_35_source_pat_all_offset;
  assign _stream_conv2d_2_source_35_source_pat_all_offset = _stream_conv2d_2_source_35_source_offset_buf + _source_stream_conv2d_2_source_35_pat_cur_offset_0 + _source_stream_conv2d_2_source_35_pat_cur_offset_1 + _source_stream_conv2d_2_source_35_pat_cur_offset_2 + _source_stream_conv2d_2_source_35_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_36_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_36_pat_stride_buf_3;
  wire _set_flag_244;
  assign _set_flag_244 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id8_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_36_source_ram_renable && (_stream_conv2d_2_source_36_source_sel == 17))? _stream_conv2d_2_source_36_source_ram_raddr : 'hx;
  assign ram_w32_l128_id8_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_36_source_ram_renable && (_stream_conv2d_2_source_36_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_245 = 1;
  wire [_tmp_245-1:0] _tmp_246;
  assign _tmp_246 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_36_source_ram_renable && (_stream_conv2d_2_source_36_source_sel == 17);
  reg [_tmp_245-1:0] __tmp_246_1;
  assign _stream_conv2d_2_source_36_source_ram_rdata = (_stream_conv2d_2_source_36_source_sel == 17)? ram_w32_l128_id8_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_554;
  assign stream_conv2d_2_source_36_data = __variable_wdata_554;
  reg [32-1:0] _stream_conv2d_2_source_36_source_pat_fsm_16;
  localparam _stream_conv2d_2_source_36_source_pat_fsm_16_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_36_source_pat_all_offset;
  assign _stream_conv2d_2_source_36_source_pat_all_offset = _stream_conv2d_2_source_36_source_offset_buf + _source_stream_conv2d_2_source_36_pat_cur_offset_0 + _source_stream_conv2d_2_source_36_pat_cur_offset_1 + _source_stream_conv2d_2_source_36_pat_cur_offset_2 + _source_stream_conv2d_2_source_36_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_2_source_37_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_2_source_37_pat_stride_buf_3;
  wire _set_flag_247;
  assign _set_flag_247 = conv2d_2_comp_fsm == 3;
  assign ram_w32_l128_id9_0_addr = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_37_source_ram_renable && (_stream_conv2d_2_source_37_source_sel == 18))? _stream_conv2d_2_source_37_source_ram_raddr : 'hx;
  assign ram_w32_l128_id9_0_enable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_37_source_ram_renable && (_stream_conv2d_2_source_37_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_248 = 1;
  wire [_tmp_248-1:0] _tmp_249;
  assign _tmp_249 = _stream_conv2d_2_stream_oready && _stream_conv2d_2_source_37_source_ram_renable && (_stream_conv2d_2_source_37_source_sel == 18);
  reg [_tmp_248-1:0] __tmp_249_1;
  assign _stream_conv2d_2_source_37_source_ram_rdata = (_stream_conv2d_2_source_37_source_sel == 18)? ram_w32_l128_id9_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_555;
  assign stream_conv2d_2_source_37_data = __variable_wdata_555;
  reg [32-1:0] _stream_conv2d_2_source_37_source_pat_fsm_17;
  localparam _stream_conv2d_2_source_37_source_pat_fsm_17_init = 0;
  wire [32-1:0] _stream_conv2d_2_source_37_source_pat_all_offset;
  assign _stream_conv2d_2_source_37_source_pat_all_offset = _stream_conv2d_2_source_37_source_offset_buf + _source_stream_conv2d_2_source_37_pat_cur_offset_0 + _source_stream_conv2d_2_source_37_pat_cur_offset_1 + _source_stream_conv2d_2_source_37_pat_cur_offset_2 + _source_stream_conv2d_2_source_37_pat_cur_offset_3;
  wire _set_flag_250;
  assign _set_flag_250 = conv2d_2_comp_fsm == 3;
  reg _tmp_251;
  reg _tmp_252;
  reg _tmp_253;
  reg _tmp_254;
  reg _tmp_255;
  reg _tmp_256;
  reg _tmp_257;
  reg _tmp_258;
  reg _tmp_259;
  reg _tmp_260;
  reg _tmp_261;
  reg _tmp_262;
  reg _tmp_263;
  reg _tmp_264;
  reg _tmp_265;
  reg _tmp_266;
  reg _tmp_267;
  reg _tmp_268;
  reg _tmp_269;
  reg _tmp_270;
  reg _tmp_271;
  reg _tmp_272;
  reg _tmp_273;
  reg _tmp_274;
  reg _tmp_275;
  reg _tmp_276;
  reg _tmp_277;
  reg _tmp_278;
  reg _tmp_279;
  reg _tmp_280;
  reg _tmp_281;
  localparam _tmp_282 = 33;
  wire [_tmp_282-1:0] _tmp_283;
  assign _tmp_283 = conv2d_2_stream_out_local + conv2d_2_out_page_comp_offset_buf;
  reg [_tmp_282-1:0] _tmp_284;
  reg [_tmp_282-1:0] _tmp_285;
  reg [_tmp_282-1:0] _tmp_286;
  reg [_tmp_282-1:0] _tmp_287;
  reg [_tmp_282-1:0] _tmp_288;
  reg [_tmp_282-1:0] _tmp_289;
  reg [_tmp_282-1:0] _tmp_290;
  reg [_tmp_282-1:0] _tmp_291;
  reg [_tmp_282-1:0] _tmp_292;
  reg [_tmp_282-1:0] _tmp_293;
  reg [_tmp_282-1:0] _tmp_294;
  reg [_tmp_282-1:0] _tmp_295;
  reg [_tmp_282-1:0] _tmp_296;
  reg [_tmp_282-1:0] _tmp_297;
  reg [_tmp_282-1:0] _tmp_298;
  reg [_tmp_282-1:0] _tmp_299;
  reg [_tmp_282-1:0] _tmp_300;
  reg [_tmp_282-1:0] _tmp_301;
  reg [_tmp_282-1:0] _tmp_302;
  reg [_tmp_282-1:0] _tmp_303;
  reg [_tmp_282-1:0] _tmp_304;
  reg [_tmp_282-1:0] _tmp_305;
  reg [_tmp_282-1:0] _tmp_306;
  reg [_tmp_282-1:0] _tmp_307;
  reg [_tmp_282-1:0] _tmp_308;
  reg [_tmp_282-1:0] _tmp_309;
  reg [_tmp_282-1:0] _tmp_310;
  reg [_tmp_282-1:0] _tmp_311;
  reg [_tmp_282-1:0] _tmp_312;
  reg [_tmp_282-1:0] _tmp_313;
  reg [_tmp_282-1:0] _tmp_314;
  reg [32-1:0] _tmp_315;
  reg [32-1:0] _tmp_316;
  reg [32-1:0] _tmp_317;
  reg [32-1:0] _tmp_318;
  reg [32-1:0] _tmp_319;
  reg [32-1:0] _tmp_320;
  reg [32-1:0] _tmp_321;
  reg [32-1:0] _tmp_322;
  reg [32-1:0] _tmp_323;
  reg [32-1:0] _tmp_324;
  reg [32-1:0] _tmp_325;
  reg [32-1:0] _tmp_326;
  reg [32-1:0] _tmp_327;
  reg [32-1:0] _tmp_328;
  reg [32-1:0] _tmp_329;
  reg [32-1:0] _tmp_330;
  reg [32-1:0] _tmp_331;
  reg [32-1:0] _tmp_332;
  reg [32-1:0] _tmp_333;
  reg [32-1:0] _tmp_334;
  reg [32-1:0] _tmp_335;
  reg [32-1:0] _tmp_336;
  reg [32-1:0] _tmp_337;
  reg [32-1:0] _tmp_338;
  reg [32-1:0] _tmp_339;
  reg [32-1:0] _tmp_340;
  reg [32-1:0] _tmp_341;
  reg [32-1:0] _tmp_342;
  reg [32-1:0] _tmp_343;
  reg [32-1:0] _tmp_344;
  reg [32-1:0] _tmp_345;
  assign ram_w32_l128_id0_0_wdata = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_sink_50_sink_wenable && (_stream_conv2d_2_sink_50_sink_sel == 19))? _stream_conv2d_2_sink_50_sink_wdata : 'hx;
  assign ram_w32_l128_id0_0_wenable = (_stream_conv2d_2_stream_oready && _stream_conv2d_2_sink_50_sink_wenable && (_stream_conv2d_2_sink_50_sink_sel == 19))? 1'd1 : 0;
  reg [32-1:0] _stream_conv2d_2_sink_50_sink_fsm_18;
  localparam _stream_conv2d_2_sink_50_sink_fsm_18_init = 0;
  wire _set_flag_346;
  assign _set_flag_346 = conv2d_2_comp_fsm == 4;
  assign _stream_conv2d_2_run_flag = (_set_flag_346)? 1 : 0;
  reg _tmp_347;
  reg _tmp_348;
  reg _tmp_349;
  assign _mul_3_source_stop = _mul_3_stream_oready && 1'd0;
  reg _tmp_350;
  reg _tmp_351;
  reg _tmp_352;
  reg _tmp_353;
  reg _tmp_354;
  reg _tmp_355;
  reg _tmp_356;
  reg _tmp_357;
  reg _tmp_358;
  reg _tmp_359;
  assign _mul_3_sink_start = _tmp_359;
  reg _tmp_360;
  reg _tmp_361;
  reg _tmp_362;
  reg _tmp_363;
  reg _tmp_364;
  reg _tmp_365;
  reg _tmp_366;
  reg _tmp_367;
  reg _tmp_368;
  reg _tmp_369;
  assign _mul_3_sink_stop = _tmp_369;
  reg _tmp_370;
  reg _tmp_371;
  reg _tmp_372;
  reg _tmp_373;
  reg _tmp_374;
  reg _tmp_375;
  reg _tmp_376;
  reg _tmp_377;
  reg _tmp_378;
  reg _tmp_379;
  assign _mul_3_sink_busy = _tmp_379;
  reg _tmp_380;
  assign _mul_3_busy = _mul_3_source_busy || _mul_3_sink_busy || _mul_3_busy_reg;
  reg _tmp_381;
  reg _tmp_382;
  reg _tmp_383;
  assign _mul_4_source_stop = _mul_4_stream_oready && 1'd0;
  reg _tmp_384;
  reg _tmp_385;
  reg _tmp_386;
  reg _tmp_387;
  reg _tmp_388;
  reg _tmp_389;
  reg _tmp_390;
  reg _tmp_391;
  reg _tmp_392;
  reg _tmp_393;
  assign _mul_4_sink_start = _tmp_393;
  reg _tmp_394;
  reg _tmp_395;
  reg _tmp_396;
  reg _tmp_397;
  reg _tmp_398;
  reg _tmp_399;
  reg _tmp_400;
  reg _tmp_401;
  reg _tmp_402;
  reg _tmp_403;
  assign _mul_4_sink_stop = _tmp_403;
  reg _tmp_404;
  reg _tmp_405;
  reg _tmp_406;
  reg _tmp_407;
  reg _tmp_408;
  reg _tmp_409;
  reg _tmp_410;
  reg _tmp_411;
  reg _tmp_412;
  reg _tmp_413;
  assign _mul_4_sink_busy = _tmp_413;
  reg _tmp_414;
  assign _mul_4_busy = _mul_4_source_busy || _mul_4_sink_busy || _mul_4_busy_reg;
  reg _tmp_415;
  reg _tmp_416;
  reg _tmp_417;
  assign _mul_5_source_stop = _mul_5_stream_oready && 1'd0;
  reg _tmp_418;
  reg _tmp_419;
  reg _tmp_420;
  reg _tmp_421;
  reg _tmp_422;
  reg _tmp_423;
  reg _tmp_424;
  reg _tmp_425;
  reg _tmp_426;
  reg _tmp_427;
  assign _mul_5_sink_start = _tmp_427;
  reg _tmp_428;
  reg _tmp_429;
  reg _tmp_430;
  reg _tmp_431;
  reg _tmp_432;
  reg _tmp_433;
  reg _tmp_434;
  reg _tmp_435;
  reg _tmp_436;
  reg _tmp_437;
  assign _mul_5_sink_stop = _tmp_437;
  reg _tmp_438;
  reg _tmp_439;
  reg _tmp_440;
  reg _tmp_441;
  reg _tmp_442;
  reg _tmp_443;
  reg _tmp_444;
  reg _tmp_445;
  reg _tmp_446;
  reg _tmp_447;
  assign _mul_5_sink_busy = _tmp_447;
  reg _tmp_448;
  assign _mul_5_busy = _mul_5_source_busy || _mul_5_sink_busy || _mul_5_busy_reg;
  reg _tmp_449;
  reg _tmp_450;
  reg _tmp_451;
  assign _mul_6_source_stop = _mul_6_stream_oready && 1'd0;
  reg _tmp_452;
  reg _tmp_453;
  reg _tmp_454;
  reg _tmp_455;
  reg _tmp_456;
  reg _tmp_457;
  reg _tmp_458;
  reg _tmp_459;
  reg _tmp_460;
  reg _tmp_461;
  assign _mul_6_sink_start = _tmp_461;
  reg _tmp_462;
  reg _tmp_463;
  reg _tmp_464;
  reg _tmp_465;
  reg _tmp_466;
  reg _tmp_467;
  reg _tmp_468;
  reg _tmp_469;
  reg _tmp_470;
  reg _tmp_471;
  assign _mul_6_sink_stop = _tmp_471;
  reg _tmp_472;
  reg _tmp_473;
  reg _tmp_474;
  reg _tmp_475;
  reg _tmp_476;
  reg _tmp_477;
  reg _tmp_478;
  reg _tmp_479;
  reg _tmp_480;
  reg _tmp_481;
  assign _mul_6_sink_busy = _tmp_481;
  reg _tmp_482;
  assign _mul_6_busy = _mul_6_source_busy || _mul_6_sink_busy || _mul_6_busy_reg;
  reg _tmp_483;
  reg _tmp_484;
  reg _tmp_485;
  assign _mul_7_source_stop = _mul_7_stream_oready && 1'd0;
  reg _tmp_486;
  reg _tmp_487;
  reg _tmp_488;
  reg _tmp_489;
  reg _tmp_490;
  reg _tmp_491;
  reg _tmp_492;
  reg _tmp_493;
  reg _tmp_494;
  reg _tmp_495;
  assign _mul_7_sink_start = _tmp_495;
  reg _tmp_496;
  reg _tmp_497;
  reg _tmp_498;
  reg _tmp_499;
  reg _tmp_500;
  reg _tmp_501;
  reg _tmp_502;
  reg _tmp_503;
  reg _tmp_504;
  reg _tmp_505;
  assign _mul_7_sink_stop = _tmp_505;
  reg _tmp_506;
  reg _tmp_507;
  reg _tmp_508;
  reg _tmp_509;
  reg _tmp_510;
  reg _tmp_511;
  reg _tmp_512;
  reg _tmp_513;
  reg _tmp_514;
  reg _tmp_515;
  assign _mul_7_sink_busy = _tmp_515;
  reg _tmp_516;
  assign _mul_7_busy = _mul_7_source_busy || _mul_7_sink_busy || _mul_7_busy_reg;
  reg _tmp_517;
  reg _tmp_518;
  reg _tmp_519;
  assign _mul_8_source_stop = _mul_8_stream_oready && 1'd0;
  reg _tmp_520;
  reg _tmp_521;
  reg _tmp_522;
  reg _tmp_523;
  reg _tmp_524;
  reg _tmp_525;
  reg _tmp_526;
  reg _tmp_527;
  reg _tmp_528;
  reg _tmp_529;
  assign _mul_8_sink_start = _tmp_529;
  reg _tmp_530;
  reg _tmp_531;
  reg _tmp_532;
  reg _tmp_533;
  reg _tmp_534;
  reg _tmp_535;
  reg _tmp_536;
  reg _tmp_537;
  reg _tmp_538;
  reg _tmp_539;
  assign _mul_8_sink_stop = _tmp_539;
  reg _tmp_540;
  reg _tmp_541;
  reg _tmp_542;
  reg _tmp_543;
  reg _tmp_544;
  reg _tmp_545;
  reg _tmp_546;
  reg _tmp_547;
  reg _tmp_548;
  reg _tmp_549;
  assign _mul_8_sink_busy = _tmp_549;
  reg _tmp_550;
  assign _mul_8_busy = _mul_8_source_busy || _mul_8_sink_busy || _mul_8_busy_reg;
  reg _tmp_551;
  reg _tmp_552;
  reg _tmp_553;
  assign _mul_9_source_stop = _mul_9_stream_oready && 1'd0;
  reg _tmp_554;
  reg _tmp_555;
  reg _tmp_556;
  reg _tmp_557;
  reg _tmp_558;
  reg _tmp_559;
  reg _tmp_560;
  reg _tmp_561;
  reg _tmp_562;
  reg _tmp_563;
  assign _mul_9_sink_start = _tmp_563;
  reg _tmp_564;
  reg _tmp_565;
  reg _tmp_566;
  reg _tmp_567;
  reg _tmp_568;
  reg _tmp_569;
  reg _tmp_570;
  reg _tmp_571;
  reg _tmp_572;
  reg _tmp_573;
  assign _mul_9_sink_stop = _tmp_573;
  reg _tmp_574;
  reg _tmp_575;
  reg _tmp_576;
  reg _tmp_577;
  reg _tmp_578;
  reg _tmp_579;
  reg _tmp_580;
  reg _tmp_581;
  reg _tmp_582;
  reg _tmp_583;
  assign _mul_9_sink_busy = _tmp_583;
  reg _tmp_584;
  assign _mul_9_busy = _mul_9_source_busy || _mul_9_sink_busy || _mul_9_busy_reg;
  reg _tmp_585;
  reg _tmp_586;
  reg _tmp_587;
  assign _mul_10_source_stop = _mul_10_stream_oready && 1'd0;
  reg _tmp_588;
  reg _tmp_589;
  reg _tmp_590;
  reg _tmp_591;
  reg _tmp_592;
  reg _tmp_593;
  reg _tmp_594;
  reg _tmp_595;
  reg _tmp_596;
  reg _tmp_597;
  assign _mul_10_sink_start = _tmp_597;
  reg _tmp_598;
  reg _tmp_599;
  reg _tmp_600;
  reg _tmp_601;
  reg _tmp_602;
  reg _tmp_603;
  reg _tmp_604;
  reg _tmp_605;
  reg _tmp_606;
  reg _tmp_607;
  assign _mul_10_sink_stop = _tmp_607;
  reg _tmp_608;
  reg _tmp_609;
  reg _tmp_610;
  reg _tmp_611;
  reg _tmp_612;
  reg _tmp_613;
  reg _tmp_614;
  reg _tmp_615;
  reg _tmp_616;
  reg _tmp_617;
  assign _mul_10_sink_busy = _tmp_617;
  reg _tmp_618;
  assign _mul_10_busy = _mul_10_source_busy || _mul_10_sink_busy || _mul_10_busy_reg;
  reg _tmp_619;
  reg _tmp_620;
  reg _tmp_621;
  assign _mul_11_source_stop = _mul_11_stream_oready && 1'd0;
  reg _tmp_622;
  reg _tmp_623;
  reg _tmp_624;
  reg _tmp_625;
  reg _tmp_626;
  reg _tmp_627;
  reg _tmp_628;
  reg _tmp_629;
  reg _tmp_630;
  reg _tmp_631;
  assign _mul_11_sink_start = _tmp_631;
  reg _tmp_632;
  reg _tmp_633;
  reg _tmp_634;
  reg _tmp_635;
  reg _tmp_636;
  reg _tmp_637;
  reg _tmp_638;
  reg _tmp_639;
  reg _tmp_640;
  reg _tmp_641;
  assign _mul_11_sink_stop = _tmp_641;
  reg _tmp_642;
  reg _tmp_643;
  reg _tmp_644;
  reg _tmp_645;
  reg _tmp_646;
  reg _tmp_647;
  reg _tmp_648;
  reg _tmp_649;
  reg _tmp_650;
  reg _tmp_651;
  assign _mul_11_sink_busy = _tmp_651;
  reg _tmp_652;
  assign _mul_11_busy = _mul_11_source_busy || _mul_11_sink_busy || _mul_11_busy_reg;
  reg _tmp_653;
  reg _tmp_654;
  reg _tmp_655;
  assign _add_tree_1_source_stop = _add_tree_1_stream_oready && 1'd0;
  reg _tmp_656;
  reg _tmp_657;
  reg _tmp_658;
  reg _tmp_659;
  assign _add_tree_1_sink_start = _tmp_659;
  reg _tmp_660;
  reg _tmp_661;
  reg _tmp_662;
  reg _tmp_663;
  assign _add_tree_1_sink_stop = _tmp_663;
  reg _tmp_664;
  reg _tmp_665;
  reg _tmp_666;
  reg _tmp_667;
  assign _add_tree_1_sink_busy = _tmp_667;
  reg _tmp_668;
  assign _add_tree_1_busy = _add_tree_1_source_busy || _add_tree_1_sink_busy || _add_tree_1_busy_reg;
  reg _tmp_669;
  reg _tmp_670;
  reg _tmp_671;
  reg _tmp_672;
  reg _tmp_673;
  reg _tmp_674;
  reg _tmp_675;
  reg _tmp_676;
  reg _tmp_677;
  reg _tmp_678;
  assign _acc_0_source_stop = _acc_0_stream_oready && 1'd0;
  reg _tmp_679;
  reg _tmp_680;
  reg _tmp_681;
  reg _tmp_682;
  reg _tmp_683;
  reg _tmp_684;
  reg _tmp_685;
  assign _acc_0_sink_start = _tmp_685;
  reg _tmp_686;
  reg _tmp_687;
  reg _tmp_688;
  reg _tmp_689;
  reg _tmp_690;
  reg _tmp_691;
  reg _tmp_692;
  assign _acc_0_sink_stop = _tmp_692;
  reg _tmp_693;
  reg _tmp_694;
  reg _tmp_695;
  reg _tmp_696;
  reg _tmp_697;
  reg _tmp_698;
  reg _tmp_699;
  assign _acc_0_sink_busy = _tmp_699;
  reg _tmp_700;
  assign _acc_0_busy = _acc_0_source_busy || _acc_0_sink_busy || _acc_0_busy_reg;
  reg _tmp_701;
  reg _tmp_702;
  reg _tmp_703;
  assign _mul_rshift_round_clip_2_source_stop = _mul_rshift_round_clip_2_stream_oready && 1'd0;
  reg _tmp_704;
  reg _tmp_705;
  reg _tmp_706;
  reg _tmp_707;
  reg _tmp_708;
  reg _tmp_709;
  reg _tmp_710;
  reg _tmp_711;
  reg _tmp_712;
  reg _tmp_713;
  assign _mul_rshift_round_clip_2_sink_start = _tmp_713;
  reg _tmp_714;
  reg _tmp_715;
  reg _tmp_716;
  reg _tmp_717;
  reg _tmp_718;
  reg _tmp_719;
  reg _tmp_720;
  reg _tmp_721;
  reg _tmp_722;
  reg _tmp_723;
  assign _mul_rshift_round_clip_2_sink_stop = _tmp_723;
  reg _tmp_724;
  reg _tmp_725;
  reg _tmp_726;
  reg _tmp_727;
  reg _tmp_728;
  reg _tmp_729;
  reg _tmp_730;
  reg _tmp_731;
  reg _tmp_732;
  reg _tmp_733;
  assign _mul_rshift_round_clip_2_sink_busy = _tmp_733;
  reg _tmp_734;
  assign _mul_rshift_round_clip_2_busy = _mul_rshift_round_clip_2_source_busy || _mul_rshift_round_clip_2_sink_busy || _mul_rshift_round_clip_2_busy_reg;
  reg _tmp_735;
  reg _tmp_736;
  reg _tmp_737;
  reg _tmp_738;
  reg _tmp_739;
  reg _tmp_740;
  reg [1-1:0] __variable_wdata_264;
  assign stream_conv2d_2__reduce_reset_data = __variable_wdata_264;
  reg _tmp_741;
  reg _tmp_742;
  reg _tmp_743;
  reg _tmp_744;
  assign _stream_conv2d_2_source_stop = _stream_conv2d_2_stream_oready && (_stream_conv2d_2_source_11_idle && _stream_conv2d_2_source_13_idle && _stream_conv2d_2_source_15_idle && _stream_conv2d_2_source_20_idle && _stream_conv2d_2_source_21_idle && _stream_conv2d_2_source_22_idle && _stream_conv2d_2_source_23_idle && _stream_conv2d_2_source_24_idle && _stream_conv2d_2_source_25_idle && _stream_conv2d_2_source_26_idle && _stream_conv2d_2_source_27_idle && _stream_conv2d_2_source_28_idle && _stream_conv2d_2_source_29_idle && _stream_conv2d_2_source_30_idle && _stream_conv2d_2_source_31_idle && _stream_conv2d_2_source_32_idle && _stream_conv2d_2_source_33_idle && _stream_conv2d_2_source_34_idle && _stream_conv2d_2_source_35_idle && _stream_conv2d_2_source_36_idle && _stream_conv2d_2_source_37_idle && _stream_conv2d_2_source_7_idle && _stream_conv2d_2_source_9_idle && (_stream_conv2d_2_fsm == 3));
  localparam _tmp_745 = 1;
  wire [_tmp_745-1:0] _tmp_746;
  assign _tmp_746 = _stream_conv2d_2_source_11_idle && _stream_conv2d_2_source_13_idle && _stream_conv2d_2_source_15_idle && _stream_conv2d_2_source_20_idle && _stream_conv2d_2_source_21_idle && _stream_conv2d_2_source_22_idle && _stream_conv2d_2_source_23_idle && _stream_conv2d_2_source_24_idle && _stream_conv2d_2_source_25_idle && _stream_conv2d_2_source_26_idle && _stream_conv2d_2_source_27_idle && _stream_conv2d_2_source_28_idle && _stream_conv2d_2_source_29_idle && _stream_conv2d_2_source_30_idle && _stream_conv2d_2_source_31_idle && _stream_conv2d_2_source_32_idle && _stream_conv2d_2_source_33_idle && _stream_conv2d_2_source_34_idle && _stream_conv2d_2_source_35_idle && _stream_conv2d_2_source_36_idle && _stream_conv2d_2_source_37_idle && _stream_conv2d_2_source_7_idle && _stream_conv2d_2_source_9_idle && (_stream_conv2d_2_fsm == 3);
  reg [_tmp_745-1:0] _tmp_747;
  localparam _tmp_748 = 1;
  wire [_tmp_748-1:0] _tmp_749;
  assign _tmp_749 = _stream_conv2d_2_source_11_idle && _stream_conv2d_2_source_13_idle && _stream_conv2d_2_source_15_idle && _stream_conv2d_2_source_20_idle && _stream_conv2d_2_source_21_idle && _stream_conv2d_2_source_22_idle && _stream_conv2d_2_source_23_idle && _stream_conv2d_2_source_24_idle && _stream_conv2d_2_source_25_idle && _stream_conv2d_2_source_26_idle && _stream_conv2d_2_source_27_idle && _stream_conv2d_2_source_28_idle && _stream_conv2d_2_source_29_idle && _stream_conv2d_2_source_30_idle && _stream_conv2d_2_source_31_idle && _stream_conv2d_2_source_32_idle && _stream_conv2d_2_source_33_idle && _stream_conv2d_2_source_34_idle && _stream_conv2d_2_source_35_idle && _stream_conv2d_2_source_36_idle && _stream_conv2d_2_source_37_idle && _stream_conv2d_2_source_7_idle && _stream_conv2d_2_source_9_idle && (_stream_conv2d_2_fsm == 3);
  reg [_tmp_748-1:0] _tmp_750;
  reg _tmp_751;
  reg _tmp_752;
  reg _tmp_753;
  reg _tmp_754;
  reg _tmp_755;
  reg _tmp_756;
  reg _tmp_757;
  reg _tmp_758;
  reg _tmp_759;
  reg _tmp_760;
  reg _tmp_761;
  reg _tmp_762;
  reg _tmp_763;
  reg _tmp_764;
  reg _tmp_765;
  reg _tmp_766;
  reg _tmp_767;
  reg _tmp_768;
  reg _tmp_769;
  reg _tmp_770;
  reg _tmp_771;
  reg _tmp_772;
  reg _tmp_773;
  reg _tmp_774;
  reg _tmp_775;
  reg _tmp_776;
  reg _tmp_777;
  reg _tmp_778;
  reg _tmp_779;
  reg _tmp_780;
  reg _tmp_781;
  assign _stream_conv2d_2_sink_start = _tmp_781;
  reg _tmp_782;
  reg _tmp_783;
  reg _tmp_784;
  reg _tmp_785;
  reg _tmp_786;
  reg _tmp_787;
  reg _tmp_788;
  reg _tmp_789;
  reg _tmp_790;
  reg _tmp_791;
  reg _tmp_792;
  reg _tmp_793;
  reg _tmp_794;
  reg _tmp_795;
  reg _tmp_796;
  reg _tmp_797;
  reg _tmp_798;
  reg _tmp_799;
  reg _tmp_800;
  reg _tmp_801;
  reg _tmp_802;
  reg _tmp_803;
  reg _tmp_804;
  reg _tmp_805;
  reg _tmp_806;
  reg _tmp_807;
  reg _tmp_808;
  reg _tmp_809;
  reg _tmp_810;
  reg _tmp_811;
  reg _tmp_812;
  assign _stream_conv2d_2_sink_stop = _tmp_812;
  reg _tmp_813;
  reg _tmp_814;
  reg _tmp_815;
  reg _tmp_816;
  reg _tmp_817;
  reg _tmp_818;
  reg _tmp_819;
  reg _tmp_820;
  reg _tmp_821;
  reg _tmp_822;
  reg _tmp_823;
  reg _tmp_824;
  reg _tmp_825;
  reg _tmp_826;
  reg _tmp_827;
  reg _tmp_828;
  reg _tmp_829;
  reg _tmp_830;
  reg _tmp_831;
  reg _tmp_832;
  reg _tmp_833;
  reg _tmp_834;
  reg _tmp_835;
  reg _tmp_836;
  reg _tmp_837;
  reg _tmp_838;
  reg _tmp_839;
  reg _tmp_840;
  reg _tmp_841;
  reg _tmp_842;
  reg _tmp_843;
  assign _stream_conv2d_2_sink_busy = _tmp_843;
  reg _tmp_844;
  assign _stream_conv2d_2_busy = _stream_conv2d_2_source_busy || _stream_conv2d_2_sink_busy || _stream_conv2d_2_busy_reg;
  wire conv2d_2_dma_out_mask_0;
  assign conv2d_2_dma_out_mask_0 = conv2d_2_out_row_count + 0 >= cparam_conv2d_2_out_num_row;
  wire [32-1:0] mask_addr_shifted_845;
  assign mask_addr_shifted_845 = conv2d_2_objaddr + (conv2d_2_out_base_offset + cparam_conv2d_2_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_846;
  assign mask_addr_masked_846 = mask_addr_shifted_845 << 2;
  reg [32-1:0] _maxi_write_req_fsm;
  localparam _maxi_write_req_fsm_init = 0;
  reg [33-1:0] _maxi_write_cur_global_size;
  reg _maxi_write_cont;
  wire [8-1:0] pack_write_req_op_sel_847;
  wire [32-1:0] pack_write_req_local_addr_848;
  wire [32-1:0] pack_write_req_local_stride_849;
  wire [33-1:0] pack_write_req_size_850;
  wire [32-1:0] pack_write_req_local_blocksize_851;
  assign pack_write_req_op_sel_847 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_848 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_849 = _maxi_write_local_stride;
  assign pack_write_req_size_850 = _maxi_write_local_size;
  assign pack_write_req_local_blocksize_851 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_852;
  assign pack_write_req_packed_852 = { pack_write_req_op_sel_847, pack_write_req_local_addr_848, pack_write_req_local_stride_849, pack_write_req_size_850, pack_write_req_local_blocksize_851 };
  localparam _tmp_853 = 1;
  wire [_tmp_853-1:0] _tmp_854;
  assign _tmp_854 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_853-1:0] __tmp_854_1;
  wire [32-1:0] mask_addr_shifted_855;
  assign mask_addr_shifted_855 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_856;
  assign mask_addr_masked_856 = mask_addr_shifted_855 << 2;
  wire [32-1:0] mask_addr_shifted_857;
  assign mask_addr_shifted_857 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_858;
  assign mask_addr_masked_858 = mask_addr_shifted_857 << 2;
  wire [32-1:0] mask_addr_shifted_859;
  assign mask_addr_shifted_859 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_860;
  assign mask_addr_masked_860 = mask_addr_shifted_859 << 2;
  wire [32-1:0] mask_addr_shifted_861;
  assign mask_addr_shifted_861 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_862;
  assign mask_addr_masked_862 = mask_addr_shifted_861 << 2;
  wire [32-1:0] mask_addr_shifted_863;
  assign mask_addr_shifted_863 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_864;
  assign mask_addr_masked_864 = mask_addr_shifted_863 << 2;
  wire [32-1:0] mask_addr_shifted_865;
  assign mask_addr_shifted_865 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_866;
  assign mask_addr_masked_866 = mask_addr_shifted_865 << 2;
  wire [8-1:0] pack_write_req_op_sel_867;
  wire [32-1:0] pack_write_req_local_addr_868;
  wire [32-1:0] pack_write_req_local_stride_869;
  wire [33-1:0] pack_write_req_size_870;
  wire [32-1:0] pack_write_req_local_blocksize_871;
  assign pack_write_req_op_sel_867 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_868 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_869 = _maxi_write_local_stride;
  assign pack_write_req_size_870 = _maxi_write_cur_global_size;
  assign pack_write_req_local_blocksize_871 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_872;
  assign pack_write_req_packed_872 = { pack_write_req_op_sel_867, pack_write_req_local_addr_868, pack_write_req_local_stride_869, pack_write_req_size_870, pack_write_req_local_blocksize_871 };
  assign _maxi_write_req_fifo_wdata = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6))? pack_write_req_packed_872 : 
                                      ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? pack_write_req_packed_852 : 'hx;
  assign _maxi_write_req_fifo_enq = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6))? (_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6) && !_maxi_write_req_fifo_almost_full : 
                                    ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? (_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full && !_maxi_write_req_fifo_almost_full : 0;
  localparam _tmp_873 = 1;
  wire [_tmp_873-1:0] _tmp_874;
  assign _tmp_874 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_873-1:0] __tmp_874_1;
  reg _maxi_cond_1_1;
  reg [32-1:0] _maxi_write_data_fsm;
  localparam _maxi_write_data_fsm_init = 0;
  reg [32-1:0] read_burst_fsm_22;
  localparam read_burst_fsm_22_init = 0;
  reg [7-1:0] read_burst_addr_875;
  reg [7-1:0] read_burst_stride_876;
  reg [33-1:0] read_burst_length_877;
  reg read_burst_rvalid_878;
  reg read_burst_rlast_879;
  localparam _tmp_880 = 1;
  wire [_tmp_880-1:0] _tmp_881;
  assign _tmp_881 = (read_burst_fsm_22 == 1) && (!read_burst_rvalid_878 || (maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0));
  reg [_tmp_880-1:0] __tmp_881_1;
  wire [32-1:0] read_burst_rdata_882;
  assign read_burst_rdata_882 = ram_w32_l128_id0_1_rdata;
  reg _maxi_cond_2_1;
  wire conv2d_2_update_filter;
  assign conv2d_2_update_filter = (cparam_conv2d_2_data_stationary == 0) && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) || (cparam_conv2d_2_data_stationary == 1) && !cparam_conv2d_2_keep_filter;
  wire conv2d_2_update_act;
  assign conv2d_2_update_act = (cparam_conv2d_2_data_stationary == 1) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count) || (cparam_conv2d_2_data_stationary == 0);
  wire conv2d_2_mux_next_dma_flag_0;
  assign conv2d_2_mux_next_dma_flag_0 = (conv2d_2_row_select == 0)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_0 : 
                                        (conv2d_2_row_select == 1)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_2 : 
                                        (conv2d_2_row_select == 2)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_1 : 1'd0;
  wire conv2d_2_mux_next_dma_flag_1;
  assign conv2d_2_mux_next_dma_flag_1 = (conv2d_2_row_select == 0)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_1 : 
                                        (conv2d_2_row_select == 1)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_0 : 
                                        (conv2d_2_row_select == 2)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_2 : 1'd0;
  wire conv2d_2_mux_next_dma_flag_2;
  assign conv2d_2_mux_next_dma_flag_2 = (conv2d_2_row_select == 0)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_2 : 
                                        (conv2d_2_row_select == 1)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_1 : 
                                        (conv2d_2_row_select == 2)? (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)? 1 : cparam_conv2d_2_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] celu_3_objaddr;
  reg [32-1:0] celu_3_arg_objaddr_0;
  reg [32-1:0] control_celu_3;
  localparam control_celu_3_init = 0;
  reg _control_celu_3_called;
  reg [32-1:0] celu_3_out_gaddr;
  reg [33-1:0] celu_3_comp_count;
  reg [32-1:0] celu_3_arg_gaddr_offset_0_0;
  reg [32-1:0] celu_3_arg_gaddr_offset_0_1;
  reg [32-1:0] celu_3_arg_gaddr_offset_0_2;
  reg [32-1:0] celu_3_arg_gaddr_offset_0_3;
  wire [32-1:0] celu_3_arg_gaddr_0;
  assign celu_3_arg_gaddr_0 = celu_3_arg_gaddr_offset_0_0 + celu_3_arg_gaddr_offset_0_1 + celu_3_arg_gaddr_offset_0_2 + celu_3_arg_gaddr_offset_0_3;
  reg [33-1:0] celu_3_arg_trip_count_0_0;
  reg [33-1:0] celu_3_arg_trip_count_0_1;
  reg [33-1:0] celu_3_arg_trip_count_0_2;
  reg [33-1:0] celu_3_arg_trip_count_0_3;
  reg [33-1:0] celu_3_arg_repeat_count_0_0;
  reg [33-1:0] celu_3_arg_repeat_count_0_1;
  reg [33-1:0] celu_3_arg_repeat_count_0_2;
  reg [33-1:0] celu_3_arg_repeat_count_0_3;
  reg celu_3_out_page;
  reg [32-1:0] celu_3_out_page_comp_offset;
  reg [32-1:0] celu_3_out_page_dma_offset;
  reg celu_3_arg_page_0;
  reg [32-1:0] celu_3_arg_page_comp_offset_0;
  reg [32-1:0] celu_3_arg_page_dma_offset_0;
  reg celu_3_skip_read;
  reg celu_3_skip_comp;
  reg celu_3_skip_write;
  wire [32-1:0] mask_addr_shifted_883;
  assign mask_addr_shifted_883 = celu_3_arg_objaddr_0 + celu_3_arg_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_884;
  assign mask_addr_masked_884 = mask_addr_shifted_883 << 2;
  assign _maxi_read_req_fifo_deq = ((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) && !_maxi_read_req_fifo_empty)? 1 : 0;
  reg [32-1:0] write_burst_fsm_23;
  localparam write_burst_fsm_23_init = 0;
  reg [7-1:0] write_burst_addr_885;
  reg [7-1:0] write_burst_stride_886;
  reg [33-1:0] write_burst_length_887;
  reg write_burst_done_888;
  assign ram_w32_l128_id0_1_addr = ((write_burst_fsm_23 == 1) && maxi_rvalid)? write_burst_addr_885 : 
                                   ((read_burst_fsm_22 == 1) && (!read_burst_rvalid_878 || (maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)))? read_burst_addr_875 : 'hx;
  assign ram_w32_l128_id0_1_wdata = ((write_burst_fsm_23 == 1) && maxi_rvalid)? maxi_rdata : 'hx;
  assign ram_w32_l128_id0_1_wenable = ((write_burst_fsm_23 == 1) && maxi_rvalid)? 1'd1 : 0;
  assign ram_w32_l128_id0_1_enable = ((write_burst_fsm_23 == 1) && maxi_rvalid)? 1'd1 : 
                                     ((read_burst_fsm_22 == 1) && (!read_burst_rvalid_878 || (maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  assign maxi_rready = (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2);
  wire [32-1:0] mask_addr_shifted_889;
  assign mask_addr_shifted_889 = celu_3_arg_objaddr_0 + celu_3_arg_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_890;
  assign mask_addr_masked_890 = mask_addr_shifted_889 << 2;
  wire [1-1:0] stream_celu_3_parameter_0_data;
  wire [32-1:0] stream_celu_3_source_1_data;
  reg __stream_celu_3_stream_ivalid_1;
  reg __stream_celu_3_stream_ivalid_2;
  reg __stream_celu_3_stream_ivalid_3;
  reg __stream_celu_3_stream_ivalid_4;
  reg __stream_celu_3_stream_ivalid_5;
  reg __stream_celu_3_stream_ivalid_6;
  reg __stream_celu_3_stream_ivalid_7;
  reg __stream_celu_3_stream_ivalid_8;
  wire [32-1:0] _reinterpretcast_src_846;
  assign _reinterpretcast_src_846 = stream_celu_3_source_1_data;
  wire signed [32-1:0] _reinterpretcast_data_846;
  assign _reinterpretcast_data_846 = _reinterpretcast_src_846;
  wire signed [32-1:0] _reinterpretcast_src_847;
  assign _reinterpretcast_src_847 = cparam_celu_3_local_0_features_scale_cparam;
  wire signed [7-1:0] _reinterpretcast_data_847;
  assign _reinterpretcast_data_847 = _reinterpretcast_src_847;
  wire signed [39-1:0] _times_mul_odata_849;
  reg signed [39-1:0] _times_mul_odata_reg_849;
  wire signed [39-1:0] _times_data_849;
  assign _times_data_849 = _times_mul_odata_reg_849;
  wire _times_mul_update_849;
  assign _times_mul_update_849 = _stream_celu_3_stream_oready;

  multiplier_1
  _times_mul_849
  (
    .CLK(CLK),
    .update(_times_mul_update_849),
    .a(_reinterpretcast_data_846),
    .b(_reinterpretcast_data_847),
    .c(_times_mul_odata_849)
  );

  wire signed [32-1:0] _reinterpretcast_src_850;
  assign _reinterpretcast_src_850 = cparam_celu_3_local_0_features_shamt_cparam;
  wire [1-1:0] _reinterpretcast_data_850;
  assign _reinterpretcast_data_850 = _reinterpretcast_src_850;
  reg [1-1:0] _greatereq_data_862;
  reg [1-1:0] __delay_data_999_reinterpretcast_850;
  reg signed [32-1:0] __delay_data_1009_reinterpretcast_846;
  reg [1-1:0] __delay_data_1000__delay_999_reinterpretcast_850;
  reg [1-1:0] __delay_data_1003_greatereq_862;
  reg signed [32-1:0] __delay_data_1010__delay_1009_reinterpretcast_846;
  reg [1-1:0] __delay_data_1001__delay_1000__delay_999_reinterpretcast_850;
  reg [1-1:0] __delay_data_1004__delay_1003_greatereq_862;
  reg signed [32-1:0] __delay_data_1011__delay_1010__delay_1009_reinterpretcast_846;
  reg signed [39-1:0] _abs_data_852;
  reg [1-1:0] __delay_data_1002__delay_1001__delay_1000___reinterpretcast_850;
  reg [1-1:0] __delay_data_1005__delay_1004__delay_1003_greatereq_862;
  reg signed [32-1:0] __delay_data_1012__delay_1011__delay_1010___reinterpretcast_846;
  reg signed [39-1:0] _sra_data_853;
  reg [1-1:0] __delay_data_1006__delay_1005__delay_1004___greatereq_862;
  reg signed [32-1:0] __delay_data_1013__delay_1012__delay_1011___reinterpretcast_846;
  wire [8-1:0] _slice_data_856;
  assign _slice_data_856 = _sra_data_853[4'd7:1'd0];
  wire [8-1:0] _lut_lut_address_857;
  assign _lut_lut_address_857 = _slice_data_856;
  wire signed [32-1:0] _lut_data_857;

  _lut_LUT_ROM_857
  _lut_lut_857
  (
    .CLK(CLK),
    .addr(_lut_lut_address_857),
    .enable(_stream_celu_3_stream_oready),
    .val(_lut_data_857)
  );

  reg [1-1:0] _greaterthan_data_858;
  reg [1-1:0] __delay_data_1007__delay_1006__delay_1005___greatereq_862;
  reg signed [32-1:0] __delay_data_1014__delay_1013__delay_1012___reinterpretcast_846;
  reg signed [33-1:0] _cond_data_860;
  reg [1-1:0] __delay_data_1008__delay_1007__delay_1006___greatereq_862;
  reg signed [32-1:0] __delay_data_1015__delay_1014__delay_1013___reinterpretcast_846;
  reg signed [33-1:0] _cond_data_864;
  wire signed [33-1:0] _reinterpretcast_src_865;
  assign _reinterpretcast_src_865 = _cond_data_864;
  wire signed [32-1:0] _reinterpretcast_data_865;
  assign _reinterpretcast_data_865 = _reinterpretcast_src_865;
  wire signed [32-1:0] stream_celu_3_sink_2_data;
  assign stream_celu_3_sink_2_data = _reinterpretcast_data_865;
  wire _set_flag_891;
  assign _set_flag_891 = control_celu_3 == 13;
  reg [1-1:0] __variable_wdata_844;
  assign stream_celu_3_parameter_0_data = __variable_wdata_844;
  wire _set_flag_892;
  assign _set_flag_892 = control_celu_3 == 13;
  assign ram_w32_l128_id0_0_addr = (_stream_celu_3_stream_oready && _stream_celu_3_source_1_source_ram_renable && (_stream_celu_3_source_1_source_sel == 1))? _stream_celu_3_source_1_source_ram_raddr : 
                                   (_stream_conv2d_2_stream_oready && _stream_conv2d_2_sink_50_sink_wenable && (_stream_conv2d_2_sink_50_sink_sel == 19))? _stream_conv2d_2_sink_50_sink_waddr : 'hx;
  assign ram_w32_l128_id0_0_enable = (_stream_celu_3_stream_oready && _stream_celu_3_source_1_source_ram_renable && (_stream_celu_3_source_1_source_sel == 1))? 1'd1 : 
                                     (_stream_conv2d_2_stream_oready && _stream_conv2d_2_sink_50_sink_wenable && (_stream_conv2d_2_sink_50_sink_sel == 19))? 1'd1 : 0;
  localparam _tmp_893 = 1;
  wire [_tmp_893-1:0] _tmp_894;
  assign _tmp_894 = _stream_celu_3_stream_oready && _stream_celu_3_source_1_source_ram_renable && (_stream_celu_3_source_1_source_sel == 1);
  reg [_tmp_893-1:0] __tmp_894_1;
  assign _stream_celu_3_source_1_source_ram_rdata = (_stream_celu_3_source_1_source_sel == 1)? ram_w32_l128_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_845;
  assign stream_celu_3_source_1_data = __variable_wdata_845;
  reg [32-1:0] _stream_celu_3_source_1_source_fsm_0;
  localparam _stream_celu_3_source_1_source_fsm_0_init = 0;
  wire _set_flag_895;
  assign _set_flag_895 = control_celu_3 == 13;
  reg _tmp_896;
  reg _tmp_897;
  reg _tmp_898;
  reg _tmp_899;
  reg _tmp_900;
  reg _tmp_901;
  reg _tmp_902;
  reg _tmp_903;
  reg _tmp_904;
  reg _tmp_905;
  reg [32-1:0] _tmp_906;
  reg [32-1:0] _tmp_907;
  reg [32-1:0] _tmp_908;
  reg [32-1:0] _tmp_909;
  reg [32-1:0] _tmp_910;
  reg [32-1:0] _tmp_911;
  reg [32-1:0] _tmp_912;
  reg [32-1:0] _tmp_913;
  reg [32-1:0] _tmp_914;
  reg [32-1:0] _tmp_915;
  reg [3-1:0] _tmp_916;
  reg [3-1:0] _tmp_917;
  reg [3-1:0] _tmp_918;
  reg [3-1:0] _tmp_919;
  reg [3-1:0] _tmp_920;
  reg [3-1:0] _tmp_921;
  reg [3-1:0] _tmp_922;
  reg [3-1:0] _tmp_923;
  reg [3-1:0] _tmp_924;
  reg [3-1:0] _tmp_925;
  assign ram_w32_l128_id1_0_addr = (_stream_celu_3_stream_oready && _stream_celu_3_sink_2_sink_wenable && (_stream_celu_3_sink_2_sink_sel == 2))? _stream_celu_3_sink_2_sink_waddr : 
                                   (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_29_source_ram_renable && (_stream_conv2d_2_source_29_source_sel == 10))? _stream_conv2d_2_source_29_source_ram_raddr : 'hx;
  assign ram_w32_l128_id1_0_wdata = (_stream_celu_3_stream_oready && _stream_celu_3_sink_2_sink_wenable && (_stream_celu_3_sink_2_sink_sel == 2))? _stream_celu_3_sink_2_sink_wdata : 'hx;
  assign ram_w32_l128_id1_0_wenable = (_stream_celu_3_stream_oready && _stream_celu_3_sink_2_sink_wenable && (_stream_celu_3_sink_2_sink_sel == 2))? 1'd1 : 0;
  assign ram_w32_l128_id1_0_enable = (_stream_celu_3_stream_oready && _stream_celu_3_sink_2_sink_wenable && (_stream_celu_3_sink_2_sink_sel == 2))? 1'd1 : 
                                     (_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_29_source_ram_renable && (_stream_conv2d_2_source_29_source_sel == 10))? 1'd1 : 0;
  reg [32-1:0] _stream_celu_3_sink_2_sink_fsm_1;
  localparam _stream_celu_3_sink_2_sink_fsm_1_init = 0;
  wire _set_flag_926;
  assign _set_flag_926 = control_celu_3 == 15;
  assign _stream_celu_3_run_flag = (_set_flag_926)? 1 : 0;
  reg _tmp_927;
  reg _tmp_928;
  reg _tmp_929;
  assign _stream_celu_3_source_stop = _stream_celu_3_stream_oready && (_stream_celu_3_source_1_idle && (_stream_celu_3_fsm == 3));
  localparam _tmp_930 = 1;
  wire [_tmp_930-1:0] _tmp_931;
  assign _tmp_931 = _stream_celu_3_source_1_idle && (_stream_celu_3_fsm == 3);
  reg [_tmp_930-1:0] _tmp_932;
  reg _tmp_933;
  reg _tmp_934;
  reg _tmp_935;
  reg _tmp_936;
  reg _tmp_937;
  reg _tmp_938;
  reg _tmp_939;
  reg _tmp_940;
  reg _tmp_941;
  reg _tmp_942;
  assign _stream_celu_3_sink_start = _tmp_942;
  reg _tmp_943;
  reg _tmp_944;
  reg _tmp_945;
  reg _tmp_946;
  reg _tmp_947;
  reg _tmp_948;
  reg _tmp_949;
  reg _tmp_950;
  reg _tmp_951;
  reg _tmp_952;
  assign _stream_celu_3_sink_stop = _tmp_952;
  reg _tmp_953;
  reg _tmp_954;
  reg _tmp_955;
  reg _tmp_956;
  reg _tmp_957;
  reg _tmp_958;
  reg _tmp_959;
  reg _tmp_960;
  reg _tmp_961;
  reg _tmp_962;
  assign _stream_celu_3_sink_busy = _tmp_962;
  reg _tmp_963;
  assign _stream_celu_3_busy = _stream_celu_3_source_busy || _stream_celu_3_sink_busy || _stream_celu_3_busy_reg;
  wire [32-1:0] mask_addr_shifted_964;
  assign mask_addr_shifted_964 = celu_3_objaddr + celu_3_out_gaddr + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_965;
  assign mask_addr_masked_965 = mask_addr_shifted_964 << 2;
  reg [32-1:0] read_burst_fsm_24;
  localparam read_burst_fsm_24_init = 0;
  reg [7-1:0] read_burst_addr_966;
  reg [7-1:0] read_burst_stride_967;
  reg [33-1:0] read_burst_length_968;
  reg read_burst_rvalid_969;
  reg read_burst_rlast_970;
  assign ram_w32_l128_id1_1_addr = ((read_burst_fsm_24 == 1) && (!read_burst_rvalid_969 || (maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)))? read_burst_addr_966 : 
                                   ((write_burst_fsm_0 == 1) && write_burst_block_ram_wvalid_47)? write_burst_addr_49 : 'hx;
  assign ram_w32_l128_id1_1_enable = ((read_burst_fsm_24 == 1) && (!read_burst_rvalid_969 || (maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                     ((write_burst_fsm_0 == 1) && write_burst_block_ram_wvalid_47)? 1'd1 : 0;
  localparam _tmp_971 = 1;
  wire [_tmp_971-1:0] _tmp_972;
  assign _tmp_972 = (read_burst_fsm_24 == 1) && (!read_burst_rvalid_969 || (maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0));
  reg [_tmp_971-1:0] __tmp_972_1;
  wire [32-1:0] read_burst_rdata_973;
  assign read_burst_rdata_973 = ram_w32_l128_id1_1_rdata;
  assign _maxi_write_req_fifo_deq = ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (_maxi_write_data_idle && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (_maxi_write_data_idle && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) && !_maxi_write_req_fifo_empty)? 1 : 0;
  reg _maxi_cond_3_1;

  always @(posedge CLK) begin
    _RESETN_inv_1 <= RESETN_inv;
    _RESETN_inv_2 <= _RESETN_inv_1;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      outstanding_wcount_0 <= 0;
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= 0;
      _maxi_read_op_sel <= 0;
      _maxi_read_global_addr <= 0;
      _maxi_read_global_size <= 0;
      _maxi_read_local_addr <= 0;
      _maxi_read_local_stride <= 0;
      _maxi_read_local_size <= 0;
      _maxi_read_local_blocksize <= 0;
      _maxi_read_req_idle <= 1;
      _maxi_read_cur_global_size <= 0;
      maxi_araddr <= 0;
      maxi_arlen <= 0;
      maxi_arvalid <= 0;
      _maxi_cond_0_1 <= 0;
      _maxi_read_data_idle <= 1;
      _maxi_read_op_sel_buf <= 0;
      _maxi_read_local_addr_buf <= 0;
      _maxi_read_local_stride_buf <= 0;
      _maxi_read_local_size_buf <= 0;
      _maxi_read_local_blocksize_buf <= 0;
      _maxi_write_op_sel <= 0;
      _maxi_write_global_addr <= 0;
      _maxi_write_global_size <= 0;
      _maxi_write_local_addr <= 0;
      _maxi_write_local_stride <= 0;
      _maxi_write_local_size <= 0;
      _maxi_write_local_blocksize <= 0;
      _maxi_write_req_idle <= 1;
      _maxi_write_cur_global_size <= 0;
      maxi_awaddr <= 0;
      maxi_awlen <= 0;
      maxi_awvalid <= 0;
      _maxi_cond_1_1 <= 0;
      _maxi_write_data_idle <= 1;
      _maxi_write_op_sel_buf <= 0;
      _maxi_write_local_addr_buf <= 0;
      _maxi_write_local_stride_buf <= 0;
      _maxi_write_size_buf <= 0;
      _maxi_write_local_blocksize_buf <= 0;
      maxi_wdata <= 0;
      maxi_wvalid <= 0;
      maxi_wlast <= 0;
      maxi_wstrb <= 0;
      _maxi_cond_2_1 <= 0;
      _maxi_cond_3_1 <= 0;
    end else begin
      if(_maxi_cond_0_1) begin
        maxi_arvalid <= 0;
      end 
      if(_maxi_cond_1_1) begin
        maxi_awvalid <= 0;
      end 
      if(_maxi_cond_2_1) begin
        maxi_wvalid <= 0;
        maxi_wlast <= 0;
      end 
      if(_maxi_cond_3_1) begin
        maxi_wvalid <= 0;
        maxi_wlast <= 0;
      end 
      if(maxi_awvalid && maxi_awready && !(maxi_bvalid && maxi_bready) && (outstanding_wcount_0 < 7)) begin
        outstanding_wcount_0 <= outstanding_wcount_0 + 1;
      end 
      if(!(maxi_awvalid && maxi_awready) && (maxi_bvalid && maxi_bready) && (outstanding_wcount_0 > 0)) begin
        outstanding_wcount_0 <= outstanding_wcount_0 - 1;
      end 
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= _saxi_register_32;
      if((control_conv2d_2 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 1;
        _maxi_read_global_addr <= mask_addr_masked_26;
        _maxi_read_global_size <= cparam_conv2d_2_filter_read_size;
        _maxi_read_local_addr <= conv2d_2_filter_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_2_filter_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_2_filter_read_block;
      end 
      if((_maxi_read_req_fsm == 0) && _maxi_read_start) begin
        _maxi_read_req_idle <= 0;
      end 
      if(_maxi_read_start && _maxi_read_req_fifo_almost_full) begin
        _maxi_read_start <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256) && ((mask_addr_masked_36 & 4095) + (_maxi_read_global_size << 2) >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_38 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_40 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256)) begin
        _maxi_read_cur_global_size <= _maxi_read_global_size;
        _maxi_read_global_size <= 0;
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && ((mask_addr_masked_42 & 4095) + 1024 >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_44 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_46 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
        _maxi_read_cur_global_size <= 256;
        _maxi_read_global_size <= _maxi_read_global_size - 256;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        maxi_araddr <= _maxi_read_global_addr;
        maxi_arlen <= _maxi_read_cur_global_size - 1;
        maxi_arvalid <= 1;
      end 
      _maxi_cond_0_1 <= 1;
      if(maxi_arvalid && !maxi_arready) begin
        maxi_arvalid <= maxi_arvalid;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        _maxi_read_global_addr <= _maxi_read_global_addr + (_maxi_read_cur_global_size << 2);
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
        _maxi_read_req_idle <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1))) begin
        _maxi_read_data_idle <= 0;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_idle <= 1;
      end 
      if((control_conv2d_2 == 10) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 2;
        _maxi_read_global_addr <= mask_addr_masked_106;
        _maxi_read_global_size <= cparam_conv2d_2_act_read_size;
        _maxi_read_local_addr <= conv2d_2_act_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_2_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_2_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2))) begin
        _maxi_read_data_idle <= 0;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_idle <= 1;
      end 
      if((control_conv2d_2 == 13) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 3;
        _maxi_read_global_addr <= mask_addr_masked_130;
        _maxi_read_global_size <= cparam_conv2d_2_act_read_size;
        _maxi_read_local_addr <= conv2d_2_act_page_dma_offset_1;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_2_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_2_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3))) begin
        _maxi_read_data_idle <= 0;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_idle <= 1;
      end 
      if((control_conv2d_2 == 16) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 4;
        _maxi_read_global_addr <= mask_addr_masked_154;
        _maxi_read_global_size <= cparam_conv2d_2_act_read_size;
        _maxi_read_local_addr <= conv2d_2_act_page_dma_offset_2;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_2_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_2_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4))) begin
        _maxi_read_data_idle <= 0;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_idle <= 1;
      end 
      if((control_conv2d_2 == 25) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_846;
        _maxi_write_global_size <= conv2d_2_next_out_write_size;
        _maxi_write_local_addr <= conv2d_2_out_laddr_offset + conv2d_2_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= conv2d_2_next_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && _maxi_write_start) begin
        _maxi_write_req_idle <= 0;
      end 
      if(_maxi_write_start && _maxi_write_req_fifo_almost_full) begin
        _maxi_write_start <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256) && ((mask_addr_masked_856 & 4095) + (_maxi_write_global_size << 2) >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_858 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_860 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256)) begin
        _maxi_write_cur_global_size <= _maxi_write_global_size;
        _maxi_write_global_size <= 0;
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && ((mask_addr_masked_862 & 4095) + 1024 >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_864 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_866 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
        _maxi_write_cur_global_size <= 256;
        _maxi_write_global_size <= _maxi_write_global_size - 256;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (outstanding_wcount_0 < 6) && ((outstanding_wcount_0 < 6) && (maxi_awready || !maxi_awvalid))) begin
        maxi_awaddr <= _maxi_write_global_addr;
        maxi_awlen <= _maxi_write_cur_global_size - 1;
        maxi_awvalid <= 1;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (outstanding_wcount_0 < 6) && ((outstanding_wcount_0 < 6) && (maxi_awready || !maxi_awvalid)) && (_maxi_write_cur_global_size == 0)) begin
        maxi_awvalid <= 0;
      end 
      _maxi_cond_1_1 <= 1;
      if(maxi_awvalid && !maxi_awready) begin
        maxi_awvalid <= maxi_awvalid;
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6))) begin
        _maxi_write_global_addr <= _maxi_write_global_addr + (_maxi_write_cur_global_size << 2);
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6)) && (_maxi_write_global_size == 0)) begin
        _maxi_write_req_idle <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (_maxi_write_data_idle && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1))) begin
        _maxi_write_data_idle <= 0;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_878 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)) && (maxi_wready || !maxi_wvalid)) begin
        maxi_wdata <= read_burst_rdata_882;
        maxi_wvalid <= 1;
        maxi_wlast <= read_burst_rlast_879 || (_maxi_write_size_buf == 1);
        maxi_wstrb <= { 4{ 1'd1 } };
      end 
      _maxi_cond_2_1 <= 1;
      if(maxi_wvalid && !maxi_wready) begin
        maxi_wvalid <= maxi_wvalid;
        maxi_wlast <= maxi_wlast;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_878 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_878 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) && read_burst_rlast_879) begin
        _maxi_write_data_idle <= 1;
      end 
      if((control_celu_3 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 5;
        _maxi_read_global_addr <= mask_addr_masked_884;
        _maxi_read_global_size <= cparam_celu_3_dma_size;
        _maxi_read_local_addr <= celu_3_arg_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_celu_3_dma_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5))) begin
        _maxi_read_data_idle <= 0;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_idle <= 1;
      end 
      if((control_celu_3 == 9) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 5;
        _maxi_read_global_addr <= mask_addr_masked_890;
        _maxi_read_global_size <= 1;
        _maxi_read_local_addr <= celu_3_arg_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= 1;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_celu_3 == 19) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 2;
        _maxi_write_global_addr <= mask_addr_masked_965;
        _maxi_write_global_size <= cparam_celu_3_dma_size;
        _maxi_write_local_addr <= celu_3_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= cparam_celu_3_dma_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (_maxi_write_data_idle && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2))) begin
        _maxi_write_data_idle <= 0;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_969 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)) && (maxi_wready || !maxi_wvalid)) begin
        maxi_wdata <= read_burst_rdata_973;
        maxi_wvalid <= 1;
        maxi_wlast <= read_burst_rlast_970 || (_maxi_write_size_buf == 1);
        maxi_wstrb <= { 4{ 1'd1 } };
      end 
      _maxi_cond_3_1 <= 1;
      if(maxi_wvalid && !maxi_wready) begin
        maxi_wvalid <= maxi_wvalid;
        maxi_wlast <= maxi_wlast;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_969 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_969 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) && read_burst_rlast_970) begin
        _maxi_write_data_idle <= 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_read_req_fifo <= 0;
      __tmp_34_1 <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full && (_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty)) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo;
      end else if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo + 1;
      end else if(_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo - 1;
      end 
      __tmp_34_1 <= _tmp_34;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_write_req_fifo <= 0;
      __tmp_854_1 <= 0;
      __tmp_874_1 <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full && (_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty)) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo;
      end else if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo + 1;
      end else if(_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo - 1;
      end 
      __tmp_854_1 <= _tmp_854;
      __tmp_874_1 <= _tmp_874;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_bvalid <= 0;
      prev_awvalid_14 <= 0;
      prev_arvalid_15 <= 0;
      writevalid_12 <= 0;
      readvalid_13 <= 0;
      addr_11 <= 0;
      saxi_rdata <= 0;
      saxi_rvalid <= 0;
      _saxi_cond_0_1 <= 0;
      _saxi_register_0 <= 0;
      _saxi_flag_0 <= 0;
      _saxi_register_1 <= 0;
      _saxi_flag_1 <= 0;
      _saxi_register_2 <= 0;
      _saxi_flag_2 <= 0;
      _saxi_register_3 <= 0;
      _saxi_flag_3 <= 0;
      _saxi_register_4 <= 0;
      _saxi_flag_4 <= 0;
      _saxi_register_5 <= 0;
      _saxi_flag_5 <= 0;
      _saxi_register_6 <= 0;
      _saxi_flag_6 <= 0;
      _saxi_register_7 <= 0;
      _saxi_flag_7 <= 0;
      _saxi_register_8 <= 0;
      _saxi_flag_8 <= 0;
      _saxi_register_9 <= 0;
      _saxi_flag_9 <= 0;
      _saxi_register_10 <= 0;
      _saxi_flag_10 <= 0;
      _saxi_register_11 <= 0;
      _saxi_flag_11 <= 0;
      _saxi_register_12 <= 0;
      _saxi_flag_12 <= 0;
      _saxi_register_13 <= 0;
      _saxi_flag_13 <= 0;
      _saxi_register_14 <= 0;
      _saxi_flag_14 <= 0;
      _saxi_register_15 <= 0;
      _saxi_flag_15 <= 0;
      _saxi_register_16 <= 0;
      _saxi_flag_16 <= 0;
      _saxi_register_17 <= 0;
      _saxi_flag_17 <= 0;
      _saxi_register_18 <= 0;
      _saxi_flag_18 <= 0;
      _saxi_register_19 <= 0;
      _saxi_flag_19 <= 0;
      _saxi_register_20 <= 0;
      _saxi_flag_20 <= 0;
      _saxi_register_21 <= 0;
      _saxi_flag_21 <= 0;
      _saxi_register_22 <= 0;
      _saxi_flag_22 <= 0;
      _saxi_register_23 <= 0;
      _saxi_flag_23 <= 0;
      _saxi_register_24 <= 0;
      _saxi_flag_24 <= 0;
      _saxi_register_25 <= 0;
      _saxi_flag_25 <= 0;
      _saxi_register_26 <= 0;
      _saxi_flag_26 <= 0;
      _saxi_register_27 <= 0;
      _saxi_flag_27 <= 0;
      _saxi_register_28 <= 0;
      _saxi_flag_28 <= 0;
      _saxi_register_29 <= 0;
      _saxi_flag_29 <= 0;
      _saxi_register_30 <= 0;
      _saxi_flag_30 <= 0;
      _saxi_register_31 <= 9600;
      _saxi_flag_31 <= 0;
      _saxi_register_32 <= 0;
      _saxi_flag_32 <= 0;
      _saxi_register_33 <= 8192;
      _saxi_flag_33 <= 0;
      _saxi_register_34 <= 0;
      _saxi_flag_34 <= 0;
      _saxi_register_35 <= 1408;
      _saxi_flag_35 <= 0;
      _saxi_register_36 <= 4352;
      _saxi_flag_36 <= 0;
      _saxi_register_11[0] <= (0 >> 0) & 1'd1;
      _saxi_register_9[0] <= (0 >> 0) & 1'd1;
      _saxi_register_11[1] <= (0 >> 1) & 1'd1;
      _saxi_register_9[1] <= (0 >> 1) & 1'd1;
      _saxi_register_11[2] <= (0 >> 2) & 1'd1;
      _saxi_register_9[2] <= (0 >> 2) & 1'd1;
      _saxi_register_11[3] <= (0 >> 3) & 1'd1;
      _saxi_register_9[3] <= (0 >> 3) & 1'd1;
      _saxi_register_11[4] <= (0 >> 4) & 1'd1;
      _saxi_register_9[4] <= (0 >> 4) & 1'd1;
      _saxi_register_11[5] <= (0 >> 5) & 1'd1;
      _saxi_register_9[5] <= (0 >> 5) & 1'd1;
      _saxi_register_11[6] <= (0 >> 6) & 1'd1;
      _saxi_register_9[6] <= (0 >> 6) & 1'd1;
      _saxi_register_11[7] <= (0 >> 7) & 1'd1;
      _saxi_register_9[7] <= (0 >> 7) & 1'd1;
      _saxi_register_11[8] <= (0 >> 8) & 1'd1;
      _saxi_register_9[8] <= (0 >> 8) & 1'd1;
      _saxi_register_11[9] <= (0 >> 9) & 1'd1;
      _saxi_register_9[9] <= (0 >> 9) & 1'd1;
      _saxi_register_11[10] <= (0 >> 10) & 1'd1;
      _saxi_register_9[10] <= (0 >> 10) & 1'd1;
      _saxi_register_11[11] <= (0 >> 11) & 1'd1;
      _saxi_register_9[11] <= (0 >> 11) & 1'd1;
      _saxi_register_11[12] <= (0 >> 12) & 1'd1;
      _saxi_register_9[12] <= (0 >> 12) & 1'd1;
      _saxi_register_11[13] <= (0 >> 13) & 1'd1;
      _saxi_register_9[13] <= (0 >> 13) & 1'd1;
      _saxi_register_11[14] <= (0 >> 14) & 1'd1;
      _saxi_register_9[14] <= (0 >> 14) & 1'd1;
      _saxi_register_11[15] <= (0 >> 15) & 1'd1;
      _saxi_register_9[15] <= (0 >> 15) & 1'd1;
      _saxi_register_11[16] <= (0 >> 16) & 1'd1;
      _saxi_register_9[16] <= (0 >> 16) & 1'd1;
      _saxi_register_11[17] <= (0 >> 17) & 1'd1;
      _saxi_register_9[17] <= (0 >> 17) & 1'd1;
      _saxi_register_11[18] <= (0 >> 18) & 1'd1;
      _saxi_register_9[18] <= (0 >> 18) & 1'd1;
      _saxi_register_11[19] <= (0 >> 19) & 1'd1;
      _saxi_register_9[19] <= (0 >> 19) & 1'd1;
      _saxi_register_11[20] <= (0 >> 20) & 1'd1;
      _saxi_register_9[20] <= (0 >> 20) & 1'd1;
      _saxi_register_11[21] <= (0 >> 21) & 1'd1;
      _saxi_register_9[21] <= (0 >> 21) & 1'd1;
      _saxi_register_11[22] <= (0 >> 22) & 1'd1;
      _saxi_register_9[22] <= (0 >> 22) & 1'd1;
      _saxi_register_11[23] <= (0 >> 23) & 1'd1;
      _saxi_register_9[23] <= (0 >> 23) & 1'd1;
      _saxi_register_11[24] <= (0 >> 24) & 1'd1;
      _saxi_register_9[24] <= (0 >> 24) & 1'd1;
      _saxi_register_11[25] <= (0 >> 25) & 1'd1;
      _saxi_register_9[25] <= (0 >> 25) & 1'd1;
      _saxi_register_11[26] <= (0 >> 26) & 1'd1;
      _saxi_register_9[26] <= (0 >> 26) & 1'd1;
      _saxi_register_11[27] <= (0 >> 27) & 1'd1;
      _saxi_register_9[27] <= (0 >> 27) & 1'd1;
      _saxi_register_11[28] <= (0 >> 28) & 1'd1;
      _saxi_register_9[28] <= (0 >> 28) & 1'd1;
      _saxi_register_11[29] <= (0 >> 29) & 1'd1;
      _saxi_register_9[29] <= (0 >> 29) & 1'd1;
      _saxi_register_11[30] <= (0 >> 30) & 1'd1;
      _saxi_register_9[30] <= (0 >> 30) & 1'd1;
      _saxi_register_11[31] <= (0 >> 31) & 1'd1;
      _saxi_register_9[31] <= (0 >> 31) & 1'd1;
      internal_state_counter <= 0;
    end else begin
      if(_saxi_cond_0_1) begin
        saxi_rvalid <= 0;
      end 
      if(saxi_bvalid && saxi_bready) begin
        saxi_bvalid <= 0;
      end 
      if(saxi_wvalid && saxi_wready) begin
        saxi_bvalid <= 1;
      end 
      prev_awvalid_14 <= saxi_awvalid;
      prev_arvalid_15 <= saxi_arvalid;
      writevalid_12 <= 0;
      readvalid_13 <= 0;
      if(saxi_awready && saxi_awvalid && !saxi_bvalid) begin
        addr_11 <= saxi_awaddr;
        writevalid_12 <= 1;
      end else if(saxi_arready && saxi_arvalid) begin
        addr_11 <= saxi_araddr;
        readvalid_13 <= 1;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid)) begin
        saxi_rdata <= axislite_rdata_17;
        saxi_rvalid <= 1;
      end 
      _saxi_cond_0_1 <= 1;
      if(saxi_rvalid && !saxi_rready) begin
        saxi_rvalid <= saxi_rvalid;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 0)) begin
        _saxi_register_0 <= axislite_resetval_19;
        _saxi_flag_0 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 1)) begin
        _saxi_register_1 <= axislite_resetval_19;
        _saxi_flag_1 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 2)) begin
        _saxi_register_2 <= axislite_resetval_19;
        _saxi_flag_2 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 3)) begin
        _saxi_register_3 <= axislite_resetval_19;
        _saxi_flag_3 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 4)) begin
        _saxi_register_4 <= axislite_resetval_19;
        _saxi_flag_4 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 5)) begin
        _saxi_register_5 <= axislite_resetval_19;
        _saxi_flag_5 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 6)) begin
        _saxi_register_6 <= axislite_resetval_19;
        _saxi_flag_6 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 7)) begin
        _saxi_register_7 <= axislite_resetval_19;
        _saxi_flag_7 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 8)) begin
        _saxi_register_8 <= axislite_resetval_19;
        _saxi_flag_8 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 9)) begin
        _saxi_register_9 <= axislite_resetval_19;
        _saxi_flag_9 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 10)) begin
        _saxi_register_10 <= axislite_resetval_19;
        _saxi_flag_10 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 11)) begin
        _saxi_register_11 <= axislite_resetval_19;
        _saxi_flag_11 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 12)) begin
        _saxi_register_12 <= axislite_resetval_19;
        _saxi_flag_12 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 13)) begin
        _saxi_register_13 <= axislite_resetval_19;
        _saxi_flag_13 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 14)) begin
        _saxi_register_14 <= axislite_resetval_19;
        _saxi_flag_14 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 15)) begin
        _saxi_register_15 <= axislite_resetval_19;
        _saxi_flag_15 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 16)) begin
        _saxi_register_16 <= axislite_resetval_19;
        _saxi_flag_16 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 17)) begin
        _saxi_register_17 <= axislite_resetval_19;
        _saxi_flag_17 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 18)) begin
        _saxi_register_18 <= axislite_resetval_19;
        _saxi_flag_18 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 19)) begin
        _saxi_register_19 <= axislite_resetval_19;
        _saxi_flag_19 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 20)) begin
        _saxi_register_20 <= axislite_resetval_19;
        _saxi_flag_20 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 21)) begin
        _saxi_register_21 <= axislite_resetval_19;
        _saxi_flag_21 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 22)) begin
        _saxi_register_22 <= axislite_resetval_19;
        _saxi_flag_22 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 23)) begin
        _saxi_register_23 <= axislite_resetval_19;
        _saxi_flag_23 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 24)) begin
        _saxi_register_24 <= axislite_resetval_19;
        _saxi_flag_24 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 25)) begin
        _saxi_register_25 <= axislite_resetval_19;
        _saxi_flag_25 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 26)) begin
        _saxi_register_26 <= axislite_resetval_19;
        _saxi_flag_26 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 27)) begin
        _saxi_register_27 <= axislite_resetval_19;
        _saxi_flag_27 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 28)) begin
        _saxi_register_28 <= axislite_resetval_19;
        _saxi_flag_28 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 29)) begin
        _saxi_register_29 <= axislite_resetval_19;
        _saxi_flag_29 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 30)) begin
        _saxi_register_30 <= axislite_resetval_19;
        _saxi_flag_30 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 31)) begin
        _saxi_register_31 <= axislite_resetval_19;
        _saxi_flag_31 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 32)) begin
        _saxi_register_32 <= axislite_resetval_19;
        _saxi_flag_32 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 33)) begin
        _saxi_register_33 <= axislite_resetval_19;
        _saxi_flag_33 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 34)) begin
        _saxi_register_34 <= axislite_resetval_19;
        _saxi_flag_34 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 35)) begin
        _saxi_register_35 <= axislite_resetval_19;
        _saxi_flag_35 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_18 && (axis_maskaddr_16 == 36)) begin
        _saxi_register_36 <= axislite_resetval_19;
        _saxi_flag_36 <= 0;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 0)) begin
        _saxi_register_0 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 1)) begin
        _saxi_register_1 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 2)) begin
        _saxi_register_2 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 3)) begin
        _saxi_register_3 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 4)) begin
        _saxi_register_4 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 5)) begin
        _saxi_register_5 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 6)) begin
        _saxi_register_6 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 7)) begin
        _saxi_register_7 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 8)) begin
        _saxi_register_8 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 9)) begin
        _saxi_register_9 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 10)) begin
        _saxi_register_10 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 11)) begin
        _saxi_register_11 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 12)) begin
        _saxi_register_12 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 13)) begin
        _saxi_register_13 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 14)) begin
        _saxi_register_14 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 15)) begin
        _saxi_register_15 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 16)) begin
        _saxi_register_16 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 17)) begin
        _saxi_register_17 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 18)) begin
        _saxi_register_18 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 19)) begin
        _saxi_register_19 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 20)) begin
        _saxi_register_20 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 21)) begin
        _saxi_register_21 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 22)) begin
        _saxi_register_22 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 23)) begin
        _saxi_register_23 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 24)) begin
        _saxi_register_24 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 25)) begin
        _saxi_register_25 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 26)) begin
        _saxi_register_26 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 27)) begin
        _saxi_register_27 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 28)) begin
        _saxi_register_28 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 29)) begin
        _saxi_register_29 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 30)) begin
        _saxi_register_30 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 31)) begin
        _saxi_register_31 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 32)) begin
        _saxi_register_32 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 33)) begin
        _saxi_register_33 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 34)) begin
        _saxi_register_34 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 35)) begin
        _saxi_register_35 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 2) && saxi_wvalid && (axis_maskaddr_16 == 36)) begin
        _saxi_register_36 <= saxi_wdata;
      end 
      if(_saxi_register_11[0] == 1) begin
        _saxi_register_11[0] <= 0;
        _saxi_register_9[0] <= 0;
      end 
      if(_saxi_register_11[1] == 1) begin
        _saxi_register_11[1] <= 0;
        _saxi_register_9[1] <= 0;
      end 
      if(_saxi_register_11[2] == 1) begin
        _saxi_register_11[2] <= 0;
        _saxi_register_9[2] <= 0;
      end 
      if(_saxi_register_11[3] == 1) begin
        _saxi_register_11[3] <= 0;
        _saxi_register_9[3] <= 0;
      end 
      if(_saxi_register_11[4] == 1) begin
        _saxi_register_11[4] <= 0;
        _saxi_register_9[4] <= 0;
      end 
      if(_saxi_register_11[5] == 1) begin
        _saxi_register_11[5] <= 0;
        _saxi_register_9[5] <= 0;
      end 
      if(_saxi_register_11[6] == 1) begin
        _saxi_register_11[6] <= 0;
        _saxi_register_9[6] <= 0;
      end 
      if(_saxi_register_11[7] == 1) begin
        _saxi_register_11[7] <= 0;
        _saxi_register_9[7] <= 0;
      end 
      if(_saxi_register_11[8] == 1) begin
        _saxi_register_11[8] <= 0;
        _saxi_register_9[8] <= 0;
      end 
      if(_saxi_register_11[9] == 1) begin
        _saxi_register_11[9] <= 0;
        _saxi_register_9[9] <= 0;
      end 
      if(_saxi_register_11[10] == 1) begin
        _saxi_register_11[10] <= 0;
        _saxi_register_9[10] <= 0;
      end 
      if(_saxi_register_11[11] == 1) begin
        _saxi_register_11[11] <= 0;
        _saxi_register_9[11] <= 0;
      end 
      if(_saxi_register_11[12] == 1) begin
        _saxi_register_11[12] <= 0;
        _saxi_register_9[12] <= 0;
      end 
      if(_saxi_register_11[13] == 1) begin
        _saxi_register_11[13] <= 0;
        _saxi_register_9[13] <= 0;
      end 
      if(_saxi_register_11[14] == 1) begin
        _saxi_register_11[14] <= 0;
        _saxi_register_9[14] <= 0;
      end 
      if(_saxi_register_11[15] == 1) begin
        _saxi_register_11[15] <= 0;
        _saxi_register_9[15] <= 0;
      end 
      if(_saxi_register_11[16] == 1) begin
        _saxi_register_11[16] <= 0;
        _saxi_register_9[16] <= 0;
      end 
      if(_saxi_register_11[17] == 1) begin
        _saxi_register_11[17] <= 0;
        _saxi_register_9[17] <= 0;
      end 
      if(_saxi_register_11[18] == 1) begin
        _saxi_register_11[18] <= 0;
        _saxi_register_9[18] <= 0;
      end 
      if(_saxi_register_11[19] == 1) begin
        _saxi_register_11[19] <= 0;
        _saxi_register_9[19] <= 0;
      end 
      if(_saxi_register_11[20] == 1) begin
        _saxi_register_11[20] <= 0;
        _saxi_register_9[20] <= 0;
      end 
      if(_saxi_register_11[21] == 1) begin
        _saxi_register_11[21] <= 0;
        _saxi_register_9[21] <= 0;
      end 
      if(_saxi_register_11[22] == 1) begin
        _saxi_register_11[22] <= 0;
        _saxi_register_9[22] <= 0;
      end 
      if(_saxi_register_11[23] == 1) begin
        _saxi_register_11[23] <= 0;
        _saxi_register_9[23] <= 0;
      end 
      if(_saxi_register_11[24] == 1) begin
        _saxi_register_11[24] <= 0;
        _saxi_register_9[24] <= 0;
      end 
      if(_saxi_register_11[25] == 1) begin
        _saxi_register_11[25] <= 0;
        _saxi_register_9[25] <= 0;
      end 
      if(_saxi_register_11[26] == 1) begin
        _saxi_register_11[26] <= 0;
        _saxi_register_9[26] <= 0;
      end 
      if(_saxi_register_11[27] == 1) begin
        _saxi_register_11[27] <= 0;
        _saxi_register_9[27] <= 0;
      end 
      if(_saxi_register_11[28] == 1) begin
        _saxi_register_11[28] <= 0;
        _saxi_register_9[28] <= 0;
      end 
      if(_saxi_register_11[29] == 1) begin
        _saxi_register_11[29] <= 0;
        _saxi_register_9[29] <= 0;
      end 
      if(_saxi_register_11[30] == 1) begin
        _saxi_register_11[30] <= 0;
        _saxi_register_9[30] <= 0;
      end 
      if(_saxi_register_11[31] == 1) begin
        _saxi_register_11[31] <= 0;
        _saxi_register_9[31] <= 0;
      end 
      if(irq_busy_edge_22) begin
        _saxi_register_9[0] <= irq_busy_edge_22;
      end 
      if(irq_extern_edge_24) begin
        _saxi_register_9[1] <= irq_extern_edge_24;
      end 
      if(main_fsm == 0) begin
        _saxi_register_5 <= 0;
        _saxi_register_6 <= 0;
        _saxi_register_7 <= 0;
      end 
      if(main_fsm == 1) begin
        internal_state_counter <= 0;
        _saxi_register_12 <= 0;
      end else if(main_fsm == _saxi_register_13) begin
        if(internal_state_counter == _saxi_register_14) begin
          internal_state_counter <= 0;
          _saxi_register_12 <= _saxi_register_12 + 1;
        end else begin
          internal_state_counter <= internal_state_counter + 1;
        end
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_0 <= 1;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_1 <= 1;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_2 <= 1;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_3 <= 1;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_4 <= 1;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 1) && 1) begin
        _saxi_register_5 <= 1;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_6 <= 1;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_7 <= 1;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_8 <= 1;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_9 <= 1;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_10 <= 1;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_11 <= 1;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_12 <= 1;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_13 <= 1;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_14 <= 1;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_15 <= 1;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_16 <= 1;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_17 <= 1;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_18 <= 1;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_19 <= 1;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_20 <= 1;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_21 <= 1;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_22 <= 1;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_23 <= 1;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_24 <= 1;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_25 <= 1;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_26 <= 1;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_27 <= 1;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_28 <= 1;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_29 <= 1;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_30 <= 1;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_31 <= 1;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_32 <= 1;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_33 <= 1;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_34 <= 1;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_35 <= 1;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_36 <= 1;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 2) && 1) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 19) && 1) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 19) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
    end
  end

  localparam _saxi_register_fsm_1 = 1;
  localparam _saxi_register_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _saxi_register_fsm <= _saxi_register_fsm_init;
      axis_maskaddr_16 <= 0;
    end else begin
      case(_saxi_register_fsm)
        _saxi_register_fsm_init: begin
          if(readvalid_13 || writevalid_12) begin
            axis_maskaddr_16 <= (addr_11 >> _saxi_shift) & _saxi_mask;
          end 
          if(readvalid_13) begin
            _saxi_register_fsm <= _saxi_register_fsm_1;
          end 
          if(writevalid_12) begin
            _saxi_register_fsm <= _saxi_register_fsm_2;
          end 
        end
        _saxi_register_fsm_1: begin
          if(saxi_rready || !saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
        _saxi_register_fsm_2: begin
          if(saxi_wvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    _rst_logic_1 <= rst_logic;
    _rst_logic_2 <= _rst_logic_1;
    RST <= rst_logic | _rst_logic_1 | _rst_logic_2;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq <= 0;
    end else begin
      irq <= |irq_20;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_busy_edge_21 <= 0;
    end else begin
      irq_busy_edge_21 <= irq_busy;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_extern_edge_23 <= 0;
    end else begin
      irq_extern_edge_23 <= irq_extern;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_881_1 <= 0;
      __tmp_894_1 <= 0;
    end else begin
      __tmp_881_1 <= _tmp_881;
      __tmp_894_1 <= _tmp_894;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_225_1 <= 0;
      __tmp_972_1 <= 0;
    end else begin
      __tmp_225_1 <= _tmp_225;
      __tmp_972_1 <= _tmp_972;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_228_1 <= 0;
    end else begin
      __tmp_228_1 <= _tmp_228;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_231_1 <= 0;
    end else begin
      __tmp_231_1 <= _tmp_231;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_234_1 <= 0;
    end else begin
      __tmp_234_1 <= _tmp_234;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_237_1 <= 0;
    end else begin
      __tmp_237_1 <= _tmp_237;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_240_1 <= 0;
    end else begin
      __tmp_240_1 <= _tmp_240;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_243_1 <= 0;
    end else begin
      __tmp_243_1 <= _tmp_243;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_246_1 <= 0;
    end else begin
      __tmp_246_1 <= _tmp_246;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_249_1 <= 0;
    end else begin
      __tmp_249_1 <= _tmp_249;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_198_1 <= 0;
    end else begin
      __tmp_198_1 <= _tmp_198;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_201_1 <= 0;
    end else begin
      __tmp_201_1 <= _tmp_201;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_204_1 <= 0;
    end else begin
      __tmp_204_1 <= _tmp_204;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_207_1 <= 0;
    end else begin
      __tmp_207_1 <= _tmp_207;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_210_1 <= 0;
    end else begin
      __tmp_210_1 <= _tmp_210;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_213_1 <= 0;
    end else begin
      __tmp_213_1 <= _tmp_213;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_216_1 <= 0;
    end else begin
      __tmp_216_1 <= _tmp_216;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_219_1 <= 0;
    end else begin
      __tmp_219_1 <= _tmp_219;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_222_1 <= 0;
    end else begin
      __tmp_222_1 <= _tmp_222;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_x_source_ram_renable <= 0;
      _acc_0_x_source_fifo_deq <= 0;
      _acc_0_x_idle <= 1;
      _acc_0_rshift_source_ram_renable <= 0;
      _acc_0_rshift_source_fifo_deq <= 0;
      _acc_0_rshift_idle <= 1;
      _acc_0_sum_sink_wenable <= 0;
      _acc_0_sum_sink_fifo_enq <= 0;
      _acc_0_valid_sink_wenable <= 0;
      _acc_0_valid_sink_fifo_enq <= 0;
      __acc_0_stream_ivalid_1 <= 0;
      __acc_0_stream_ivalid_2 <= 0;
      __acc_0_stream_ivalid_3 <= 0;
      __acc_0_stream_ivalid_4 <= 0;
      __acc_0_stream_ivalid_5 <= 0;
      _greaterthan_data_3 <= 0;
      _minus_data_5 <= 0;
      _reduceadd_data_16 <= 1'sd0;
      _reduceadd_count_16 <= 0;
      _reduceadd_prev_count_max_16 <= 0;
      _pulse_data_18 <= 1'sd0;
      _pulse_count_18 <= 0;
      _pulse_prev_count_max_18 <= 0;
      __delay_data_814__variable_1 <= 0;
      _sll_data_7 <= 0;
      __delay_data_811_greaterthan_3 <= 0;
      __delay_data_812_reduceadd_16 <= 0;
      __delay_data_815__delay_814__variable_1 <= 0;
      __delay_data_818_pulse_18 <= 0;
      _cond_data_13 <= 0;
      __delay_data_813__delay_812_reduceadd_16 <= 0;
      __delay_data_816__delay_815__delay_814__variable_1 <= 0;
      __delay_data_819__delay_818_pulse_18 <= 0;
      _plus_data_20 <= 0;
      __delay_data_817__delay_816__delay_815__delay_814__variable_1 <= 0;
      __delay_data_820__delay_819__delay_818_pulse_18 <= 0;
      _sra_data_21 <= 0;
      __delay_data_821__delay_820__delay_819__delay_818_pulse_18 <= 0;
      __variable_wdata_15 <= 0;
      __variable_wdata_0 <= 0;
      __variable_wdata_1 <= 0;
      __variable_wdata_2 <= 0;
      _tmp_669 <= 0;
      _tmp_670 <= 0;
      _tmp_671 <= 0;
      _tmp_672 <= 0;
      _tmp_673 <= 0;
      _tmp_674 <= 0;
      _tmp_675 <= 0;
      _tmp_676 <= 0;
      _tmp_677 <= 0;
      _tmp_678 <= 0;
      _tmp_679 <= 0;
      _tmp_680 <= 0;
      _tmp_681 <= 0;
      _tmp_682 <= 0;
      _tmp_683 <= 0;
      _tmp_684 <= 0;
      _tmp_685 <= 0;
      _tmp_686 <= 0;
      _tmp_687 <= 0;
      _tmp_688 <= 0;
      _tmp_689 <= 0;
      _tmp_690 <= 0;
      _tmp_691 <= 0;
      _tmp_692 <= 0;
      _tmp_693 <= 0;
      _tmp_694 <= 0;
      _tmp_695 <= 0;
      _tmp_696 <= 0;
      _tmp_697 <= 0;
      _tmp_698 <= 0;
      _tmp_699 <= 0;
      _tmp_700 <= 0;
      _acc_0_busy_reg <= 0;
    end else begin
      if(_acc_0_stream_oready) begin
        _acc_0_x_source_ram_renable <= 0;
        _acc_0_x_source_fifo_deq <= 0;
      end 
      _acc_0_x_idle <= _acc_0_x_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_rshift_source_ram_renable <= 0;
        _acc_0_rshift_source_fifo_deq <= 0;
      end 
      _acc_0_rshift_idle <= _acc_0_rshift_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_sum_sink_wenable <= 0;
        _acc_0_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        _acc_0_valid_sink_wenable <= 0;
        _acc_0_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_1 <= _acc_0_stream_ivalid;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_2 <= __acc_0_stream_ivalid_1;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_3 <= __acc_0_stream_ivalid_2;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_4 <= __acc_0_stream_ivalid_3;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_5 <= __acc_0_stream_ivalid_4;
      end 
      if(_acc_0_stream_oready) begin
        _greaterthan_data_3 <= acc_0_rshift_data > 1'sd0;
      end 
      if(_acc_0_stream_oready) begin
        _minus_data_5 <= acc_0_rshift_data - 2'sd1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _reduceadd_reset_cond_16) begin
        _reduceadd_data_16 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_count_16 <= (_reduceadd_current_count_16 >= acc_0_size_data - 1)? 0 : _reduceadd_current_count_16 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_prev_count_max_16 <= _reduceadd_current_count_16 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_data_16 <= _reduceadd_current_data_16 + acc_0_x_data;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _pulse_reset_cond_18) begin
        _pulse_data_18 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_count_18 <= (_pulse_current_count_18 >= acc_0_size_data - 1)? 0 : _pulse_current_count_18 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_prev_count_max_18 <= _pulse_current_count_18 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_data_18 <= _pulse_current_count_18 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_814__variable_1 <= acc_0_rshift_data;
      end 
      if(_acc_0_stream_oready) begin
        _sll_data_7 <= 2'sd1 << _minus_data_5;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_811_greaterthan_3 <= _greaterthan_data_3;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_812_reduceadd_16 <= _reduceadd_data_16;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_815__delay_814__variable_1 <= __delay_data_814__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_818_pulse_18 <= _pulse_data_18;
      end 
      if(_acc_0_stream_oready) begin
        _cond_data_13 <= (__delay_data_811_greaterthan_3)? _sll_data_7 : 1'sd0;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_813__delay_812_reduceadd_16 <= __delay_data_812_reduceadd_16;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_816__delay_815__delay_814__variable_1 <= __delay_data_815__delay_814__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_819__delay_818_pulse_18 <= __delay_data_818_pulse_18;
      end 
      if(_acc_0_stream_oready) begin
        _plus_data_20 <= __delay_data_813__delay_812_reduceadd_16 + _cond_data_13;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_817__delay_816__delay_815__delay_814__variable_1 <= __delay_data_816__delay_815__delay_814__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_820__delay_819__delay_818_pulse_18 <= __delay_data_819__delay_818_pulse_18;
      end 
      if(_acc_0_stream_oready) begin
        _sra_data_21 <= _plus_data_20 >>> __delay_data_817__delay_816__delay_815__delay_814__variable_1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_821__delay_820__delay_819__delay_818_pulse_18 <= __delay_data_820__delay_819__delay_818_pulse_18;
      end 
      if(__stream_conv2d_2_stream_ivalid_13 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_15 <= __delay_data_905__delay_904__delay_903____variable_264;
      end 
      if(__stream_conv2d_2_stream_ivalid_13 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_0 <= __substreamoutput_data_809;
      end 
      if(__stream_conv2d_2_stream_ivalid_13 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_1 <= __delay_data_917__delay_916__delay_915__delay_914___plus_822;
      end 
      if(__stream_conv2d_2_stream_ivalid_13 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_2 <= __delay_data_930__delay_929__delay_928____variable_259;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_669 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_670 <= _tmp_669;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_671 <= _tmp_670;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_672 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_673 <= _tmp_672;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_674 <= _tmp_673;
      end 
      if(_acc_0_stream_oready && _tmp_674) begin
        __variable_wdata_15 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_675 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_676 <= _tmp_675;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_677 <= _tmp_676;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_678 <= _tmp_677;
      end 
      if(_acc_0_stream_oready && _tmp_678) begin
        __variable_wdata_15 <= 0;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        __variable_wdata_15 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_679 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_680 <= _tmp_679;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_681 <= _tmp_680;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_682 <= _tmp_681;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_683 <= _tmp_682;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_684 <= _tmp_683;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_685 <= _tmp_684;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_686 <= _acc_0_source_stop;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_687 <= _tmp_686;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_688 <= _tmp_687;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_689 <= _tmp_688;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_690 <= _tmp_689;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_691 <= _tmp_690;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_692 <= _tmp_691;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_693 <= _acc_0_source_busy;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_694 <= _tmp_693;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_695 <= _tmp_694;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_696 <= _tmp_695;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_697 <= _tmp_696;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_698 <= _tmp_697;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_699 <= _tmp_698;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_700 <= _acc_0_sink_busy;
      end 
      if(!_acc_0_sink_busy && _tmp_700) begin
        _acc_0_busy_reg <= 0;
      end 
      if(_acc_0_source_busy) begin
        _acc_0_busy_reg <= 1;
      end 
    end
  end

  localparam _acc_0_fsm_1 = 1;
  localparam _acc_0_fsm_2 = 2;
  localparam _acc_0_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_fsm <= _acc_0_fsm_init;
      _acc_0_source_start <= 0;
      _acc_0_source_busy <= 0;
      _acc_0_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_13 && _stream_conv2d_2_stream_oready) begin
        _acc_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _acc_0_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_acc_0_stream_oready && _tmp_671) begin
        _acc_0_stream_ivalid <= 1;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        _acc_0_stream_ivalid <= 0;
      end 
      case(_acc_0_fsm)
        _acc_0_fsm_init: begin
          if(_acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
        _acc_0_fsm_1: begin
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_source_start <= 0;
            _acc_0_source_busy <= 1;
          end 
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_2;
          end 
        end
        _acc_0_fsm_2: begin
          if(_acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_3;
          end 
        end
        _acc_0_fsm_3: begin
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_source_busy <= 0;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_fsm <= _acc_0_fsm_init;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_1_var0_source_ram_renable <= 0;
      _add_tree_1_var0_source_fifo_deq <= 0;
      _add_tree_1_var0_idle <= 1;
      _add_tree_1_var1_source_ram_renable <= 0;
      _add_tree_1_var1_source_fifo_deq <= 0;
      _add_tree_1_var1_idle <= 1;
      _add_tree_1_var2_source_ram_renable <= 0;
      _add_tree_1_var2_source_fifo_deq <= 0;
      _add_tree_1_var2_idle <= 1;
      _add_tree_1_var3_source_ram_renable <= 0;
      _add_tree_1_var3_source_fifo_deq <= 0;
      _add_tree_1_var3_idle <= 1;
      _add_tree_1_var4_source_ram_renable <= 0;
      _add_tree_1_var4_source_fifo_deq <= 0;
      _add_tree_1_var4_idle <= 1;
      _add_tree_1_var5_source_ram_renable <= 0;
      _add_tree_1_var5_source_fifo_deq <= 0;
      _add_tree_1_var5_idle <= 1;
      _add_tree_1_var6_source_ram_renable <= 0;
      _add_tree_1_var6_source_fifo_deq <= 0;
      _add_tree_1_var6_idle <= 1;
      _add_tree_1_var7_source_ram_renable <= 0;
      _add_tree_1_var7_source_fifo_deq <= 0;
      _add_tree_1_var7_idle <= 1;
      _add_tree_1_var8_source_ram_renable <= 0;
      _add_tree_1_var8_source_fifo_deq <= 0;
      _add_tree_1_var8_idle <= 1;
      _add_tree_1_sum_sink_wenable <= 0;
      _add_tree_1_sum_sink_fifo_enq <= 0;
      __add_tree_1_stream_ivalid_1 <= 0;
      __add_tree_1_stream_ivalid_2 <= 0;
      __plusn_data_32 <= 0;
      __plusn_data_33 <= 0;
      __plusn_data_34 <= 0;
      __plusn_data_35 <= 0;
      __variable_wdata_22 <= 0;
      __variable_wdata_23 <= 0;
      __variable_wdata_24 <= 0;
      __variable_wdata_25 <= 0;
      __variable_wdata_26 <= 0;
      __variable_wdata_27 <= 0;
      __variable_wdata_28 <= 0;
      __variable_wdata_29 <= 0;
      __variable_wdata_30 <= 0;
      _tmp_653 <= 0;
      _tmp_654 <= 0;
      _tmp_655 <= 0;
      _tmp_656 <= 0;
      _tmp_657 <= 0;
      _tmp_658 <= 0;
      _tmp_659 <= 0;
      _tmp_660 <= 0;
      _tmp_661 <= 0;
      _tmp_662 <= 0;
      _tmp_663 <= 0;
      _tmp_664 <= 0;
      _tmp_665 <= 0;
      _tmp_666 <= 0;
      _tmp_667 <= 0;
      _tmp_668 <= 0;
      _add_tree_1_busy_reg <= 0;
    end else begin
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var0_source_ram_renable <= 0;
        _add_tree_1_var0_source_fifo_deq <= 0;
      end 
      _add_tree_1_var0_idle <= _add_tree_1_var0_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var1_source_ram_renable <= 0;
        _add_tree_1_var1_source_fifo_deq <= 0;
      end 
      _add_tree_1_var1_idle <= _add_tree_1_var1_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var2_source_ram_renable <= 0;
        _add_tree_1_var2_source_fifo_deq <= 0;
      end 
      _add_tree_1_var2_idle <= _add_tree_1_var2_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var3_source_ram_renable <= 0;
        _add_tree_1_var3_source_fifo_deq <= 0;
      end 
      _add_tree_1_var3_idle <= _add_tree_1_var3_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var4_source_ram_renable <= 0;
        _add_tree_1_var4_source_fifo_deq <= 0;
      end 
      _add_tree_1_var4_idle <= _add_tree_1_var4_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var5_source_ram_renable <= 0;
        _add_tree_1_var5_source_fifo_deq <= 0;
      end 
      _add_tree_1_var5_idle <= _add_tree_1_var5_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var6_source_ram_renable <= 0;
        _add_tree_1_var6_source_fifo_deq <= 0;
      end 
      _add_tree_1_var6_idle <= _add_tree_1_var6_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var7_source_ram_renable <= 0;
        _add_tree_1_var7_source_fifo_deq <= 0;
      end 
      _add_tree_1_var7_idle <= _add_tree_1_var7_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_var8_source_ram_renable <= 0;
        _add_tree_1_var8_source_fifo_deq <= 0;
      end 
      _add_tree_1_var8_idle <= _add_tree_1_var8_idle;
      if(_add_tree_1_stream_oready) begin
        _add_tree_1_sum_sink_wenable <= 0;
        _add_tree_1_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_1_stream_oready) begin
        __add_tree_1_stream_ivalid_1 <= _add_tree_1_stream_ivalid;
      end 
      if(_add_tree_1_stream_oready) begin
        __add_tree_1_stream_ivalid_2 <= __add_tree_1_stream_ivalid_1;
      end 
      if(_add_tree_1_stream_oready) begin
        __plusn_data_32 <= add_tree_1_var0_data + add_tree_1_var1_data + add_tree_1_var2_data;
      end 
      if(_add_tree_1_stream_oready) begin
        __plusn_data_33 <= add_tree_1_var3_data + add_tree_1_var4_data + add_tree_1_var5_data;
      end 
      if(_add_tree_1_stream_oready) begin
        __plusn_data_34 <= add_tree_1_var6_data + add_tree_1_var7_data + add_tree_1_var8_data;
      end 
      if(_add_tree_1_stream_oready) begin
        __plusn_data_35 <= __plusn_data_32 + __plusn_data_33 + __plusn_data_34;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_22 <= __substreamoutput_data_655;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_23 <= __substreamoutput_data_674;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_24 <= __substreamoutput_data_693;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_25 <= __substreamoutput_data_712;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_26 <= __substreamoutput_data_731;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_27 <= __substreamoutput_data_750;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_28 <= __substreamoutput_data_769;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_29 <= __substreamoutput_data_788;
      end 
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_30 <= __substreamoutput_data_807;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_653 <= _add_tree_1_source_start;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_654 <= _tmp_653;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_655 <= _tmp_654;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_656 <= _add_tree_1_source_start;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_657 <= _tmp_656;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_658 <= _tmp_657;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_659 <= _tmp_658;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_660 <= _add_tree_1_source_stop;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_661 <= _tmp_660;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_662 <= _tmp_661;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_663 <= _tmp_662;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_664 <= _add_tree_1_source_busy;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_665 <= _tmp_664;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_666 <= _tmp_665;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_667 <= _tmp_666;
      end 
      if(_add_tree_1_stream_oready) begin
        _tmp_668 <= _add_tree_1_sink_busy;
      end 
      if(!_add_tree_1_sink_busy && _tmp_668) begin
        _add_tree_1_busy_reg <= 0;
      end 
      if(_add_tree_1_source_busy) begin
        _add_tree_1_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_1_fsm_1 = 1;
  localparam _add_tree_1_fsm_2 = 2;
  localparam _add_tree_1_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_1_fsm <= _add_tree_1_fsm_init;
      _add_tree_1_source_start <= 0;
      _add_tree_1_source_busy <= 0;
      _add_tree_1_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_10 && _stream_conv2d_2_stream_oready) begin
        _add_tree_1_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _add_tree_1_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_add_tree_1_stream_oready && _tmp_655) begin
        _add_tree_1_stream_ivalid <= 1;
      end 
      if(_add_tree_1_stream_oready && 1'd0) begin
        _add_tree_1_stream_ivalid <= 0;
      end 
      case(_add_tree_1_fsm)
        _add_tree_1_fsm_init: begin
          if(_add_tree_1_run_flag) begin
            _add_tree_1_source_start <= 1;
          end 
          if(_add_tree_1_run_flag) begin
            _add_tree_1_fsm <= _add_tree_1_fsm_1;
          end 
        end
        _add_tree_1_fsm_1: begin
          if(_add_tree_1_source_start && _add_tree_1_stream_oready) begin
            _add_tree_1_source_start <= 0;
            _add_tree_1_source_busy <= 1;
          end 
          if(_add_tree_1_source_start && _add_tree_1_stream_oready) begin
            _add_tree_1_fsm <= _add_tree_1_fsm_2;
          end 
        end
        _add_tree_1_fsm_2: begin
          if(_add_tree_1_stream_oready) begin
            _add_tree_1_fsm <= _add_tree_1_fsm_3;
          end 
        end
        _add_tree_1_fsm_3: begin
          if(_add_tree_1_stream_oready && 1'd0) begin
            _add_tree_1_source_busy <= 0;
          end 
          if(_add_tree_1_stream_oready && 1'd0 && _add_tree_1_run_flag) begin
            _add_tree_1_source_start <= 1;
          end 
          if(_add_tree_1_stream_oready && 1'd0) begin
            _add_tree_1_fsm <= _add_tree_1_fsm_init;
          end 
          if(_add_tree_1_stream_oready && 1'd0 && _add_tree_1_run_flag) begin
            _add_tree_1_fsm <= _add_tree_1_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_2_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_2_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_2_x_idle <= 1;
      _mul_rshift_round_clip_2_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_2_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_2_y_idle <= 1;
      _mul_rshift_round_clip_2_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_2_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_2_rshift_idle <= 1;
      _mul_rshift_round_clip_2_z_sink_wenable <= 0;
      _mul_rshift_round_clip_2_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_2_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_39 <= 0;
      __delay_data_827_sll_45 <= 0;
      __delay_data_831__variable_38 <= 0;
      __delay_data_835_eq_57 <= 0;
      __delay_data_828__delay_827_sll_45 <= 0;
      __delay_data_832__delay_831__variable_38 <= 0;
      __delay_data_836__delay_835_eq_57 <= 0;
      __delay_data_829__delay_828__delay_827_sll_45 <= 0;
      __delay_data_833__delay_832__delay_831__variable_38 <= 0;
      __delay_data_837__delay_836__delay_835_eq_57 <= 0;
      __delay_data_830__delay_829__delay_828__delay_827_sll_45 <= 0;
      __delay_data_834__delay_833__delay_832__delay_831__variable_38 <= 0;
      __delay_data_838__delay_837__delay_836__delay_835_eq_57 <= 0;
      _cond_data_58 <= 0;
      _greaterthan_data_59 <= 0;
      _lessthan_data_63 <= 0;
      _greatereq_data_67 <= 0;
      __delay_data_839_cond_58 <= 0;
      _cond_data_61 <= 0;
      _cond_data_65 <= 0;
      __delay_data_840_greatereq_67 <= 0;
      _cond_data_69 <= 0;
      __variable_wdata_36 <= 0;
      __variable_wdata_37 <= 0;
      __variable_wdata_38 <= 0;
      _tmp_701 <= 0;
      _tmp_702 <= 0;
      _tmp_703 <= 0;
      _tmp_704 <= 0;
      _tmp_705 <= 0;
      _tmp_706 <= 0;
      _tmp_707 <= 0;
      _tmp_708 <= 0;
      _tmp_709 <= 0;
      _tmp_710 <= 0;
      _tmp_711 <= 0;
      _tmp_712 <= 0;
      _tmp_713 <= 0;
      _tmp_714 <= 0;
      _tmp_715 <= 0;
      _tmp_716 <= 0;
      _tmp_717 <= 0;
      _tmp_718 <= 0;
      _tmp_719 <= 0;
      _tmp_720 <= 0;
      _tmp_721 <= 0;
      _tmp_722 <= 0;
      _tmp_723 <= 0;
      _tmp_724 <= 0;
      _tmp_725 <= 0;
      _tmp_726 <= 0;
      _tmp_727 <= 0;
      _tmp_728 <= 0;
      _tmp_729 <= 0;
      _tmp_730 <= 0;
      _tmp_731 <= 0;
      _tmp_732 <= 0;
      _tmp_733 <= 0;
      _tmp_734 <= 0;
      _mul_rshift_round_clip_2_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _mul_rshift_round_clip_2_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_2_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_2_x_idle <= _mul_rshift_round_clip_2_x_idle;
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _mul_rshift_round_clip_2_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_2_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_2_y_idle <= _mul_rshift_round_clip_2_y_idle;
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _mul_rshift_round_clip_2_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_2_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_2_rshift_idle <= _mul_rshift_round_clip_2_rshift_idle;
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _mul_rshift_round_clip_2_z_sink_wenable <= 0;
        _mul_rshift_round_clip_2_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_1 <= _mul_rshift_round_clip_2_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_2 <= __mul_rshift_round_clip_2_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_3 <= __mul_rshift_round_clip_2_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_4 <= __mul_rshift_round_clip_2_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_5 <= __mul_rshift_round_clip_2_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_6 <= __mul_rshift_round_clip_2_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_7 <= __mul_rshift_round_clip_2_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __mul_rshift_round_clip_2_stream_ivalid_8 <= __mul_rshift_round_clip_2_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _times_mul_odata_reg_39 <= _times_mul_odata_39;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_827_sll_45 <= _sll_data_45;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_831__variable_38 <= mul_rshift_round_clip_2_rshift_data;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_835_eq_57 <= _eq_data_57;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_828__delay_827_sll_45 <= __delay_data_827_sll_45;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_832__delay_831__variable_38 <= __delay_data_831__variable_38;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_836__delay_835_eq_57 <= __delay_data_835_eq_57;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_829__delay_828__delay_827_sll_45 <= __delay_data_828__delay_827_sll_45;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_833__delay_832__delay_831__variable_38 <= __delay_data_832__delay_831__variable_38;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_837__delay_836__delay_835_eq_57 <= __delay_data_836__delay_835_eq_57;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_830__delay_829__delay_828__delay_827_sll_45 <= __delay_data_829__delay_828__delay_827_sll_45;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_834__delay_833__delay_832__delay_831__variable_38 <= __delay_data_833__delay_832__delay_831__variable_38;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_838__delay_837__delay_836__delay_835_eq_57 <= __delay_data_837__delay_836__delay_835_eq_57;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _cond_data_58 <= (__delay_data_838__delay_837__delay_836__delay_835_eq_57)? _times_data_39 : _sra_data_55;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _greaterthan_data_59 <= _cond_data_58 > 32'sd2147483647;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _lessthan_data_63 <= _cond_data_58 < -32'sd2147483647;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _greatereq_data_67 <= _cond_data_58 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_839_cond_58 <= _cond_data_58;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _cond_data_61 <= (_greaterthan_data_59)? 32'sd2147483647 : __delay_data_839_cond_58;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _cond_data_65 <= (_lessthan_data_63)? -32'sd2147483647 : __delay_data_839_cond_58;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        __delay_data_840_greatereq_67 <= _greatereq_data_67;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _cond_data_69 <= (__delay_data_840_greatereq_67)? _cond_data_61 : _cond_data_65;
      end 
      if(__stream_conv2d_2_stream_ivalid_20 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_36 <= _plus_data_825;
      end 
      if(__stream_conv2d_2_stream_ivalid_20 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_37 <= __delay_data_969__delay_968__delay_967__delay_966___cond_287;
      end 
      if(__stream_conv2d_2_stream_ivalid_20 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_38 <= __delay_data_988__delay_987__delay_986__delay_985___plus_841;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_701 <= _mul_rshift_round_clip_2_source_start;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_702 <= _tmp_701;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_703 <= _tmp_702;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_704 <= _mul_rshift_round_clip_2_source_start;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_705 <= _tmp_704;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_706 <= _tmp_705;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_707 <= _tmp_706;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_708 <= _tmp_707;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_709 <= _tmp_708;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_710 <= _tmp_709;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_711 <= _tmp_710;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_712 <= _tmp_711;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_713 <= _tmp_712;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_714 <= _mul_rshift_round_clip_2_source_stop;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_715 <= _tmp_714;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_716 <= _tmp_715;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_717 <= _tmp_716;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_718 <= _tmp_717;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_719 <= _tmp_718;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_720 <= _tmp_719;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_721 <= _tmp_720;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_722 <= _tmp_721;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_723 <= _tmp_722;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_724 <= _mul_rshift_round_clip_2_source_busy;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_725 <= _tmp_724;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_726 <= _tmp_725;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_727 <= _tmp_726;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_728 <= _tmp_727;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_729 <= _tmp_728;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_730 <= _tmp_729;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_731 <= _tmp_730;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_732 <= _tmp_731;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_733 <= _tmp_732;
      end 
      if(_mul_rshift_round_clip_2_stream_oready) begin
        _tmp_734 <= _mul_rshift_round_clip_2_sink_busy;
      end 
      if(!_mul_rshift_round_clip_2_sink_busy && _tmp_734) begin
        _mul_rshift_round_clip_2_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_2_source_busy) begin
        _mul_rshift_round_clip_2_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_rshift_round_clip_2_fsm_1 = 1;
  localparam _mul_rshift_round_clip_2_fsm_2 = 2;
  localparam _mul_rshift_round_clip_2_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_2_fsm <= _mul_rshift_round_clip_2_fsm_init;
      _mul_rshift_round_clip_2_source_start <= 0;
      _mul_rshift_round_clip_2_source_busy <= 0;
      _mul_rshift_round_clip_2_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_20 && _stream_conv2d_2_stream_oready) begin
        _mul_rshift_round_clip_2_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_rshift_round_clip_2_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_rshift_round_clip_2_stream_oready && _tmp_703) begin
        _mul_rshift_round_clip_2_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_2_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_2_stream_ivalid <= 0;
      end 
      case(_mul_rshift_round_clip_2_fsm)
        _mul_rshift_round_clip_2_fsm_init: begin
          if(_mul_rshift_round_clip_2_run_flag) begin
            _mul_rshift_round_clip_2_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_2_run_flag) begin
            _mul_rshift_round_clip_2_fsm <= _mul_rshift_round_clip_2_fsm_1;
          end 
        end
        _mul_rshift_round_clip_2_fsm_1: begin
          if(_mul_rshift_round_clip_2_source_start && _mul_rshift_round_clip_2_stream_oready) begin
            _mul_rshift_round_clip_2_source_start <= 0;
            _mul_rshift_round_clip_2_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_2_source_start && _mul_rshift_round_clip_2_stream_oready) begin
            _mul_rshift_round_clip_2_fsm <= _mul_rshift_round_clip_2_fsm_2;
          end 
        end
        _mul_rshift_round_clip_2_fsm_2: begin
          if(_mul_rshift_round_clip_2_stream_oready) begin
            _mul_rshift_round_clip_2_fsm <= _mul_rshift_round_clip_2_fsm_3;
          end 
        end
        _mul_rshift_round_clip_2_fsm_3: begin
          if(_mul_rshift_round_clip_2_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_2_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_2_stream_oready && 1'd0 && _mul_rshift_round_clip_2_run_flag) begin
            _mul_rshift_round_clip_2_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_2_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_2_fsm <= _mul_rshift_round_clip_2_fsm_init;
          end 
          if(_mul_rshift_round_clip_2_stream_oready && 1'd0 && _mul_rshift_round_clip_2_run_flag) begin
            _mul_rshift_round_clip_2_fsm <= _mul_rshift_round_clip_2_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_3_x_source_ram_renable <= 0;
      _mul_3_x_source_fifo_deq <= 0;
      _mul_3_x_idle <= 1;
      _mul_3_y_source_ram_renable <= 0;
      _mul_3_y_source_fifo_deq <= 0;
      _mul_3_y_idle <= 1;
      _mul_3_rshift_source_ram_renable <= 0;
      _mul_3_rshift_source_fifo_deq <= 0;
      _mul_3_rshift_idle <= 1;
      _mul_3_z_sink_wenable <= 0;
      _mul_3_z_sink_fifo_enq <= 0;
      __mul_3_stream_ivalid_1 <= 0;
      __mul_3_stream_ivalid_2 <= 0;
      __mul_3_stream_ivalid_3 <= 0;
      __mul_3_stream_ivalid_4 <= 0;
      __mul_3_stream_ivalid_5 <= 0;
      __mul_3_stream_ivalid_6 <= 0;
      __mul_3_stream_ivalid_7 <= 0;
      __mul_3_stream_ivalid_8 <= 0;
      _greaterthan_data_73 <= 0;
      _minus_data_75 <= 0;
      _greatereq_data_86 <= 0;
      __delay_data_641__variable_70 <= 0;
      __delay_data_644__variable_71 <= 0;
      __delay_data_647__variable_72 <= 0;
      _sll_data_77 <= 0;
      __delay_data_638_greaterthan_73 <= 0;
      __delay_data_639_greatereq_86 <= 0;
      __delay_data_642__delay_641__variable_70 <= 0;
      __delay_data_645__delay_644__variable_71 <= 0;
      __delay_data_648__delay_647__variable_72 <= 0;
      _cond_data_83 <= 0;
      __delay_data_640__delay_639_greatereq_86 <= 0;
      __delay_data_643__delay_642__delay_641__variable_70 <= 0;
      __delay_data_646__delay_645__delay_644__variable_71 <= 0;
      __delay_data_649__delay_648__delay_647__variable_72 <= 0;
      __muladd_madd_odata_reg_89 <= 0;
      __delay_data_650__delay_649__delay_648__delay_647__variable_72 <= 0;
      __delay_data_651__delay_650__delay_649__delay_648____variable_72 <= 0;
      __delay_data_652__delay_651__delay_650__delay_649____variable_72 <= 0;
      __delay_data_653__delay_652__delay_651__delay_650____variable_72 <= 0;
      _sra_data_90 <= 0;
      __variable_wdata_70 <= 0;
      __variable_wdata_71 <= 0;
      __variable_wdata_72 <= 0;
      _tmp_347 <= 0;
      _tmp_348 <= 0;
      _tmp_349 <= 0;
      _tmp_350 <= 0;
      _tmp_351 <= 0;
      _tmp_352 <= 0;
      _tmp_353 <= 0;
      _tmp_354 <= 0;
      _tmp_355 <= 0;
      _tmp_356 <= 0;
      _tmp_357 <= 0;
      _tmp_358 <= 0;
      _tmp_359 <= 0;
      _tmp_360 <= 0;
      _tmp_361 <= 0;
      _tmp_362 <= 0;
      _tmp_363 <= 0;
      _tmp_364 <= 0;
      _tmp_365 <= 0;
      _tmp_366 <= 0;
      _tmp_367 <= 0;
      _tmp_368 <= 0;
      _tmp_369 <= 0;
      _tmp_370 <= 0;
      _tmp_371 <= 0;
      _tmp_372 <= 0;
      _tmp_373 <= 0;
      _tmp_374 <= 0;
      _tmp_375 <= 0;
      _tmp_376 <= 0;
      _tmp_377 <= 0;
      _tmp_378 <= 0;
      _tmp_379 <= 0;
      _tmp_380 <= 0;
      _mul_3_busy_reg <= 0;
    end else begin
      if(_mul_3_stream_oready) begin
        _mul_3_x_source_ram_renable <= 0;
        _mul_3_x_source_fifo_deq <= 0;
      end 
      _mul_3_x_idle <= _mul_3_x_idle;
      if(_mul_3_stream_oready) begin
        _mul_3_y_source_ram_renable <= 0;
        _mul_3_y_source_fifo_deq <= 0;
      end 
      _mul_3_y_idle <= _mul_3_y_idle;
      if(_mul_3_stream_oready) begin
        _mul_3_rshift_source_ram_renable <= 0;
        _mul_3_rshift_source_fifo_deq <= 0;
      end 
      _mul_3_rshift_idle <= _mul_3_rshift_idle;
      if(_mul_3_stream_oready) begin
        _mul_3_z_sink_wenable <= 0;
        _mul_3_z_sink_fifo_enq <= 0;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_1 <= _mul_3_stream_ivalid;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_2 <= __mul_3_stream_ivalid_1;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_3 <= __mul_3_stream_ivalid_2;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_4 <= __mul_3_stream_ivalid_3;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_5 <= __mul_3_stream_ivalid_4;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_6 <= __mul_3_stream_ivalid_5;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_7 <= __mul_3_stream_ivalid_6;
      end 
      if(_mul_3_stream_oready) begin
        __mul_3_stream_ivalid_8 <= __mul_3_stream_ivalid_7;
      end 
      if(_mul_3_stream_oready) begin
        _greaterthan_data_73 <= mul_3_rshift_data > 1'sd0;
      end 
      if(_mul_3_stream_oready) begin
        _minus_data_75 <= mul_3_rshift_data - 2'sd1;
      end 
      if(_mul_3_stream_oready) begin
        _greatereq_data_86 <= mul_3_x_data >= 1'sd0;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_641__variable_70 <= mul_3_x_data;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_644__variable_71 <= mul_3_y_data;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_647__variable_72 <= mul_3_rshift_data;
      end 
      if(_mul_3_stream_oready) begin
        _sll_data_77 <= 2'sd1 << _minus_data_75;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_638_greaterthan_73 <= _greaterthan_data_73;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_639_greatereq_86 <= _greatereq_data_86;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_642__delay_641__variable_70 <= __delay_data_641__variable_70;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_645__delay_644__variable_71 <= __delay_data_644__variable_71;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_648__delay_647__variable_72 <= __delay_data_647__variable_72;
      end 
      if(_mul_3_stream_oready) begin
        _cond_data_83 <= (__delay_data_638_greaterthan_73)? _sll_data_77 : 1'sd0;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_640__delay_639_greatereq_86 <= __delay_data_639_greatereq_86;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_643__delay_642__delay_641__variable_70 <= __delay_data_642__delay_641__variable_70;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_646__delay_645__delay_644__variable_71 <= __delay_data_645__delay_644__variable_71;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_649__delay_648__delay_647__variable_72 <= __delay_data_648__delay_647__variable_72;
      end 
      if(_mul_3_stream_oready) begin
        __muladd_madd_odata_reg_89 <= __muladd_madd_odata_89;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_650__delay_649__delay_648__delay_647__variable_72 <= __delay_data_649__delay_648__delay_647__variable_72;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_651__delay_650__delay_649__delay_648____variable_72 <= __delay_data_650__delay_649__delay_648__delay_647__variable_72;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_652__delay_651__delay_650__delay_649____variable_72 <= __delay_data_651__delay_650__delay_649__delay_648____variable_72;
      end 
      if(_mul_3_stream_oready) begin
        __delay_data_653__delay_652__delay_651__delay_650____variable_72 <= __delay_data_652__delay_651__delay_650__delay_649____variable_72;
      end 
      if(_mul_3_stream_oready) begin
        _sra_data_90 <= __muladd_data_89 >>> __delay_data_653__delay_652__delay_651__delay_650____variable_72;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_70 <= _cond_data_620;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_71 <= __delay_data_876_reinterpretcast_592;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_72 <= _plus_data_654;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_347 <= _mul_3_source_start;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_348 <= _tmp_347;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_349 <= _tmp_348;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_350 <= _mul_3_source_start;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_351 <= _tmp_350;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_352 <= _tmp_351;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_353 <= _tmp_352;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_354 <= _tmp_353;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_355 <= _tmp_354;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_356 <= _tmp_355;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_357 <= _tmp_356;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_358 <= _tmp_357;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_359 <= _tmp_358;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_360 <= _mul_3_source_stop;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_361 <= _tmp_360;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_362 <= _tmp_361;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_363 <= _tmp_362;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_364 <= _tmp_363;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_365 <= _tmp_364;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_366 <= _tmp_365;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_367 <= _tmp_366;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_368 <= _tmp_367;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_369 <= _tmp_368;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_370 <= _mul_3_source_busy;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_371 <= _tmp_370;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_372 <= _tmp_371;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_373 <= _tmp_372;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_374 <= _tmp_373;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_375 <= _tmp_374;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_376 <= _tmp_375;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_377 <= _tmp_376;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_378 <= _tmp_377;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_379 <= _tmp_378;
      end 
      if(_mul_3_stream_oready) begin
        _tmp_380 <= _mul_3_sink_busy;
      end 
      if(!_mul_3_sink_busy && _tmp_380) begin
        _mul_3_busy_reg <= 0;
      end 
      if(_mul_3_source_busy) begin
        _mul_3_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_3_fsm_1 = 1;
  localparam _mul_3_fsm_2 = 2;
  localparam _mul_3_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_3_fsm <= _mul_3_fsm_init;
      _mul_3_source_start <= 0;
      _mul_3_source_busy <= 0;
      _mul_3_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_3_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_3_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_3_stream_oready && _tmp_349) begin
        _mul_3_stream_ivalid <= 1;
      end 
      if(_mul_3_stream_oready && 1'd0) begin
        _mul_3_stream_ivalid <= 0;
      end 
      case(_mul_3_fsm)
        _mul_3_fsm_init: begin
          if(_mul_3_run_flag) begin
            _mul_3_source_start <= 1;
          end 
          if(_mul_3_run_flag) begin
            _mul_3_fsm <= _mul_3_fsm_1;
          end 
        end
        _mul_3_fsm_1: begin
          if(_mul_3_source_start && _mul_3_stream_oready) begin
            _mul_3_source_start <= 0;
            _mul_3_source_busy <= 1;
          end 
          if(_mul_3_source_start && _mul_3_stream_oready) begin
            _mul_3_fsm <= _mul_3_fsm_2;
          end 
        end
        _mul_3_fsm_2: begin
          if(_mul_3_stream_oready) begin
            _mul_3_fsm <= _mul_3_fsm_3;
          end 
        end
        _mul_3_fsm_3: begin
          if(_mul_3_stream_oready && 1'd0) begin
            _mul_3_source_busy <= 0;
          end 
          if(_mul_3_stream_oready && 1'd0 && _mul_3_run_flag) begin
            _mul_3_source_start <= 1;
          end 
          if(_mul_3_stream_oready && 1'd0) begin
            _mul_3_fsm <= _mul_3_fsm_init;
          end 
          if(_mul_3_stream_oready && 1'd0 && _mul_3_run_flag) begin
            _mul_3_fsm <= _mul_3_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_4_x_source_ram_renable <= 0;
      _mul_4_x_source_fifo_deq <= 0;
      _mul_4_x_idle <= 1;
      _mul_4_y_source_ram_renable <= 0;
      _mul_4_y_source_fifo_deq <= 0;
      _mul_4_y_idle <= 1;
      _mul_4_rshift_source_ram_renable <= 0;
      _mul_4_rshift_source_fifo_deq <= 0;
      _mul_4_rshift_idle <= 1;
      _mul_4_z_sink_wenable <= 0;
      _mul_4_z_sink_fifo_enq <= 0;
      __mul_4_stream_ivalid_1 <= 0;
      __mul_4_stream_ivalid_2 <= 0;
      __mul_4_stream_ivalid_3 <= 0;
      __mul_4_stream_ivalid_4 <= 0;
      __mul_4_stream_ivalid_5 <= 0;
      __mul_4_stream_ivalid_6 <= 0;
      __mul_4_stream_ivalid_7 <= 0;
      __mul_4_stream_ivalid_8 <= 0;
      _greaterthan_data_94 <= 0;
      _minus_data_96 <= 0;
      _greatereq_data_107 <= 0;
      __delay_data_660__variable_91 <= 0;
      __delay_data_663__variable_92 <= 0;
      __delay_data_666__variable_93 <= 0;
      _sll_data_98 <= 0;
      __delay_data_657_greaterthan_94 <= 0;
      __delay_data_658_greatereq_107 <= 0;
      __delay_data_661__delay_660__variable_91 <= 0;
      __delay_data_664__delay_663__variable_92 <= 0;
      __delay_data_667__delay_666__variable_93 <= 0;
      _cond_data_104 <= 0;
      __delay_data_659__delay_658_greatereq_107 <= 0;
      __delay_data_662__delay_661__delay_660__variable_91 <= 0;
      __delay_data_665__delay_664__delay_663__variable_92 <= 0;
      __delay_data_668__delay_667__delay_666__variable_93 <= 0;
      __muladd_madd_odata_reg_110 <= 0;
      __delay_data_669__delay_668__delay_667__delay_666__variable_93 <= 0;
      __delay_data_670__delay_669__delay_668__delay_667____variable_93 <= 0;
      __delay_data_671__delay_670__delay_669__delay_668____variable_93 <= 0;
      __delay_data_672__delay_671__delay_670__delay_669____variable_93 <= 0;
      _sra_data_111 <= 0;
      __variable_wdata_91 <= 0;
      __variable_wdata_92 <= 0;
      __variable_wdata_93 <= 0;
      _tmp_381 <= 0;
      _tmp_382 <= 0;
      _tmp_383 <= 0;
      _tmp_384 <= 0;
      _tmp_385 <= 0;
      _tmp_386 <= 0;
      _tmp_387 <= 0;
      _tmp_388 <= 0;
      _tmp_389 <= 0;
      _tmp_390 <= 0;
      _tmp_391 <= 0;
      _tmp_392 <= 0;
      _tmp_393 <= 0;
      _tmp_394 <= 0;
      _tmp_395 <= 0;
      _tmp_396 <= 0;
      _tmp_397 <= 0;
      _tmp_398 <= 0;
      _tmp_399 <= 0;
      _tmp_400 <= 0;
      _tmp_401 <= 0;
      _tmp_402 <= 0;
      _tmp_403 <= 0;
      _tmp_404 <= 0;
      _tmp_405 <= 0;
      _tmp_406 <= 0;
      _tmp_407 <= 0;
      _tmp_408 <= 0;
      _tmp_409 <= 0;
      _tmp_410 <= 0;
      _tmp_411 <= 0;
      _tmp_412 <= 0;
      _tmp_413 <= 0;
      _tmp_414 <= 0;
      _mul_4_busy_reg <= 0;
    end else begin
      if(_mul_4_stream_oready) begin
        _mul_4_x_source_ram_renable <= 0;
        _mul_4_x_source_fifo_deq <= 0;
      end 
      _mul_4_x_idle <= _mul_4_x_idle;
      if(_mul_4_stream_oready) begin
        _mul_4_y_source_ram_renable <= 0;
        _mul_4_y_source_fifo_deq <= 0;
      end 
      _mul_4_y_idle <= _mul_4_y_idle;
      if(_mul_4_stream_oready) begin
        _mul_4_rshift_source_ram_renable <= 0;
        _mul_4_rshift_source_fifo_deq <= 0;
      end 
      _mul_4_rshift_idle <= _mul_4_rshift_idle;
      if(_mul_4_stream_oready) begin
        _mul_4_z_sink_wenable <= 0;
        _mul_4_z_sink_fifo_enq <= 0;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_1 <= _mul_4_stream_ivalid;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_2 <= __mul_4_stream_ivalid_1;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_3 <= __mul_4_stream_ivalid_2;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_4 <= __mul_4_stream_ivalid_3;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_5 <= __mul_4_stream_ivalid_4;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_6 <= __mul_4_stream_ivalid_5;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_7 <= __mul_4_stream_ivalid_6;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_8 <= __mul_4_stream_ivalid_7;
      end 
      if(_mul_4_stream_oready) begin
        _greaterthan_data_94 <= mul_4_rshift_data > 1'sd0;
      end 
      if(_mul_4_stream_oready) begin
        _minus_data_96 <= mul_4_rshift_data - 2'sd1;
      end 
      if(_mul_4_stream_oready) begin
        _greatereq_data_107 <= mul_4_x_data >= 1'sd0;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_660__variable_91 <= mul_4_x_data;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_663__variable_92 <= mul_4_y_data;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_666__variable_93 <= mul_4_rshift_data;
      end 
      if(_mul_4_stream_oready) begin
        _sll_data_98 <= 2'sd1 << _minus_data_96;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_657_greaterthan_94 <= _greaterthan_data_94;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_658_greatereq_107 <= _greatereq_data_107;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_661__delay_660__variable_91 <= __delay_data_660__variable_91;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_664__delay_663__variable_92 <= __delay_data_663__variable_92;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_667__delay_666__variable_93 <= __delay_data_666__variable_93;
      end 
      if(_mul_4_stream_oready) begin
        _cond_data_104 <= (__delay_data_657_greaterthan_94)? _sll_data_98 : 1'sd0;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_659__delay_658_greatereq_107 <= __delay_data_658_greatereq_107;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_662__delay_661__delay_660__variable_91 <= __delay_data_661__delay_660__variable_91;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_665__delay_664__delay_663__variable_92 <= __delay_data_664__delay_663__variable_92;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_668__delay_667__delay_666__variable_93 <= __delay_data_667__delay_666__variable_93;
      end 
      if(_mul_4_stream_oready) begin
        __muladd_madd_odata_reg_110 <= __muladd_madd_odata_110;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_669__delay_668__delay_667__delay_666__variable_93 <= __delay_data_668__delay_667__delay_666__variable_93;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_670__delay_669__delay_668__delay_667____variable_93 <= __delay_data_669__delay_668__delay_667__delay_666__variable_93;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_671__delay_670__delay_669__delay_668____variable_93 <= __delay_data_670__delay_669__delay_668__delay_667____variable_93;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_672__delay_671__delay_670__delay_669____variable_93 <= __delay_data_671__delay_670__delay_669__delay_668____variable_93;
      end 
      if(_mul_4_stream_oready) begin
        _sra_data_111 <= __muladd_data_110 >>> __delay_data_672__delay_671__delay_670__delay_669____variable_93;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_91 <= _cond_data_622;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_92 <= __delay_data_878_reinterpretcast_593;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_93 <= _plus_data_673;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_381 <= _mul_4_source_start;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_382 <= _tmp_381;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_383 <= _tmp_382;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_384 <= _mul_4_source_start;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_385 <= _tmp_384;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_386 <= _tmp_385;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_387 <= _tmp_386;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_388 <= _tmp_387;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_389 <= _tmp_388;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_390 <= _tmp_389;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_391 <= _tmp_390;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_392 <= _tmp_391;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_393 <= _tmp_392;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_394 <= _mul_4_source_stop;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_395 <= _tmp_394;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_396 <= _tmp_395;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_397 <= _tmp_396;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_398 <= _tmp_397;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_399 <= _tmp_398;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_400 <= _tmp_399;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_401 <= _tmp_400;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_402 <= _tmp_401;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_403 <= _tmp_402;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_404 <= _mul_4_source_busy;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_405 <= _tmp_404;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_406 <= _tmp_405;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_407 <= _tmp_406;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_408 <= _tmp_407;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_409 <= _tmp_408;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_410 <= _tmp_409;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_411 <= _tmp_410;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_412 <= _tmp_411;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_413 <= _tmp_412;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_414 <= _mul_4_sink_busy;
      end 
      if(!_mul_4_sink_busy && _tmp_414) begin
        _mul_4_busy_reg <= 0;
      end 
      if(_mul_4_source_busy) begin
        _mul_4_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_4_fsm_1 = 1;
  localparam _mul_4_fsm_2 = 2;
  localparam _mul_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_4_fsm <= _mul_4_fsm_init;
      _mul_4_source_start <= 0;
      _mul_4_source_busy <= 0;
      _mul_4_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_4_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_4_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_4_stream_oready && _tmp_383) begin
        _mul_4_stream_ivalid <= 1;
      end 
      if(_mul_4_stream_oready && 1'd0) begin
        _mul_4_stream_ivalid <= 0;
      end 
      case(_mul_4_fsm)
        _mul_4_fsm_init: begin
          if(_mul_4_run_flag) begin
            _mul_4_source_start <= 1;
          end 
          if(_mul_4_run_flag) begin
            _mul_4_fsm <= _mul_4_fsm_1;
          end 
        end
        _mul_4_fsm_1: begin
          if(_mul_4_source_start && _mul_4_stream_oready) begin
            _mul_4_source_start <= 0;
            _mul_4_source_busy <= 1;
          end 
          if(_mul_4_source_start && _mul_4_stream_oready) begin
            _mul_4_fsm <= _mul_4_fsm_2;
          end 
        end
        _mul_4_fsm_2: begin
          if(_mul_4_stream_oready) begin
            _mul_4_fsm <= _mul_4_fsm_3;
          end 
        end
        _mul_4_fsm_3: begin
          if(_mul_4_stream_oready && 1'd0) begin
            _mul_4_source_busy <= 0;
          end 
          if(_mul_4_stream_oready && 1'd0 && _mul_4_run_flag) begin
            _mul_4_source_start <= 1;
          end 
          if(_mul_4_stream_oready && 1'd0) begin
            _mul_4_fsm <= _mul_4_fsm_init;
          end 
          if(_mul_4_stream_oready && 1'd0 && _mul_4_run_flag) begin
            _mul_4_fsm <= _mul_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_x_source_ram_renable <= 0;
      _mul_5_x_source_fifo_deq <= 0;
      _mul_5_x_idle <= 1;
      _mul_5_y_source_ram_renable <= 0;
      _mul_5_y_source_fifo_deq <= 0;
      _mul_5_y_idle <= 1;
      _mul_5_rshift_source_ram_renable <= 0;
      _mul_5_rshift_source_fifo_deq <= 0;
      _mul_5_rshift_idle <= 1;
      _mul_5_z_sink_wenable <= 0;
      _mul_5_z_sink_fifo_enq <= 0;
      __mul_5_stream_ivalid_1 <= 0;
      __mul_5_stream_ivalid_2 <= 0;
      __mul_5_stream_ivalid_3 <= 0;
      __mul_5_stream_ivalid_4 <= 0;
      __mul_5_stream_ivalid_5 <= 0;
      __mul_5_stream_ivalid_6 <= 0;
      __mul_5_stream_ivalid_7 <= 0;
      __mul_5_stream_ivalid_8 <= 0;
      _greaterthan_data_115 <= 0;
      _minus_data_117 <= 0;
      _greatereq_data_128 <= 0;
      __delay_data_679__variable_112 <= 0;
      __delay_data_682__variable_113 <= 0;
      __delay_data_685__variable_114 <= 0;
      _sll_data_119 <= 0;
      __delay_data_676_greaterthan_115 <= 0;
      __delay_data_677_greatereq_128 <= 0;
      __delay_data_680__delay_679__variable_112 <= 0;
      __delay_data_683__delay_682__variable_113 <= 0;
      __delay_data_686__delay_685__variable_114 <= 0;
      _cond_data_125 <= 0;
      __delay_data_678__delay_677_greatereq_128 <= 0;
      __delay_data_681__delay_680__delay_679__variable_112 <= 0;
      __delay_data_684__delay_683__delay_682__variable_113 <= 0;
      __delay_data_687__delay_686__delay_685__variable_114 <= 0;
      __muladd_madd_odata_reg_131 <= 0;
      __delay_data_688__delay_687__delay_686____variable_114 <= 0;
      __delay_data_689__delay_688__delay_687____variable_114 <= 0;
      __delay_data_690__delay_689__delay_688____variable_114 <= 0;
      __delay_data_691__delay_690__delay_689____variable_114 <= 0;
      _sra_data_132 <= 0;
      __variable_wdata_112 <= 0;
      __variable_wdata_113 <= 0;
      __variable_wdata_114 <= 0;
      _tmp_415 <= 0;
      _tmp_416 <= 0;
      _tmp_417 <= 0;
      _tmp_418 <= 0;
      _tmp_419 <= 0;
      _tmp_420 <= 0;
      _tmp_421 <= 0;
      _tmp_422 <= 0;
      _tmp_423 <= 0;
      _tmp_424 <= 0;
      _tmp_425 <= 0;
      _tmp_426 <= 0;
      _tmp_427 <= 0;
      _tmp_428 <= 0;
      _tmp_429 <= 0;
      _tmp_430 <= 0;
      _tmp_431 <= 0;
      _tmp_432 <= 0;
      _tmp_433 <= 0;
      _tmp_434 <= 0;
      _tmp_435 <= 0;
      _tmp_436 <= 0;
      _tmp_437 <= 0;
      _tmp_438 <= 0;
      _tmp_439 <= 0;
      _tmp_440 <= 0;
      _tmp_441 <= 0;
      _tmp_442 <= 0;
      _tmp_443 <= 0;
      _tmp_444 <= 0;
      _tmp_445 <= 0;
      _tmp_446 <= 0;
      _tmp_447 <= 0;
      _tmp_448 <= 0;
      _mul_5_busy_reg <= 0;
    end else begin
      if(_mul_5_stream_oready) begin
        _mul_5_x_source_ram_renable <= 0;
        _mul_5_x_source_fifo_deq <= 0;
      end 
      _mul_5_x_idle <= _mul_5_x_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_y_source_ram_renable <= 0;
        _mul_5_y_source_fifo_deq <= 0;
      end 
      _mul_5_y_idle <= _mul_5_y_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_rshift_source_ram_renable <= 0;
        _mul_5_rshift_source_fifo_deq <= 0;
      end 
      _mul_5_rshift_idle <= _mul_5_rshift_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_z_sink_wenable <= 0;
        _mul_5_z_sink_fifo_enq <= 0;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_1 <= _mul_5_stream_ivalid;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_2 <= __mul_5_stream_ivalid_1;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_3 <= __mul_5_stream_ivalid_2;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_4 <= __mul_5_stream_ivalid_3;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_5 <= __mul_5_stream_ivalid_4;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_6 <= __mul_5_stream_ivalid_5;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_7 <= __mul_5_stream_ivalid_6;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_8 <= __mul_5_stream_ivalid_7;
      end 
      if(_mul_5_stream_oready) begin
        _greaterthan_data_115 <= mul_5_rshift_data > 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        _minus_data_117 <= mul_5_rshift_data - 2'sd1;
      end 
      if(_mul_5_stream_oready) begin
        _greatereq_data_128 <= mul_5_x_data >= 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_679__variable_112 <= mul_5_x_data;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_682__variable_113 <= mul_5_y_data;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_685__variable_114 <= mul_5_rshift_data;
      end 
      if(_mul_5_stream_oready) begin
        _sll_data_119 <= 2'sd1 << _minus_data_117;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_676_greaterthan_115 <= _greaterthan_data_115;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_677_greatereq_128 <= _greatereq_data_128;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_680__delay_679__variable_112 <= __delay_data_679__variable_112;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_683__delay_682__variable_113 <= __delay_data_682__variable_113;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_686__delay_685__variable_114 <= __delay_data_685__variable_114;
      end 
      if(_mul_5_stream_oready) begin
        _cond_data_125 <= (__delay_data_676_greaterthan_115)? _sll_data_119 : 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_678__delay_677_greatereq_128 <= __delay_data_677_greatereq_128;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_681__delay_680__delay_679__variable_112 <= __delay_data_680__delay_679__variable_112;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_684__delay_683__delay_682__variable_113 <= __delay_data_683__delay_682__variable_113;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_687__delay_686__delay_685__variable_114 <= __delay_data_686__delay_685__variable_114;
      end 
      if(_mul_5_stream_oready) begin
        __muladd_madd_odata_reg_131 <= __muladd_madd_odata_131;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_688__delay_687__delay_686____variable_114 <= __delay_data_687__delay_686__delay_685__variable_114;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_689__delay_688__delay_687____variable_114 <= __delay_data_688__delay_687__delay_686____variable_114;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_690__delay_689__delay_688____variable_114 <= __delay_data_689__delay_688__delay_687____variable_114;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_691__delay_690__delay_689____variable_114 <= __delay_data_690__delay_689__delay_688____variable_114;
      end 
      if(_mul_5_stream_oready) begin
        _sra_data_132 <= __muladd_data_131 >>> __delay_data_691__delay_690__delay_689____variable_114;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_112 <= _cond_data_624;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_113 <= __delay_data_880_reinterpretcast_594;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_114 <= _plus_data_692;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_415 <= _mul_5_source_start;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_416 <= _tmp_415;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_417 <= _tmp_416;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_418 <= _mul_5_source_start;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_419 <= _tmp_418;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_420 <= _tmp_419;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_421 <= _tmp_420;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_422 <= _tmp_421;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_423 <= _tmp_422;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_424 <= _tmp_423;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_425 <= _tmp_424;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_426 <= _tmp_425;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_427 <= _tmp_426;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_428 <= _mul_5_source_stop;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_429 <= _tmp_428;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_430 <= _tmp_429;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_431 <= _tmp_430;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_432 <= _tmp_431;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_433 <= _tmp_432;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_434 <= _tmp_433;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_435 <= _tmp_434;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_436 <= _tmp_435;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_437 <= _tmp_436;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_438 <= _mul_5_source_busy;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_439 <= _tmp_438;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_440 <= _tmp_439;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_441 <= _tmp_440;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_442 <= _tmp_441;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_443 <= _tmp_442;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_444 <= _tmp_443;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_445 <= _tmp_444;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_446 <= _tmp_445;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_447 <= _tmp_446;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_448 <= _mul_5_sink_busy;
      end 
      if(!_mul_5_sink_busy && _tmp_448) begin
        _mul_5_busy_reg <= 0;
      end 
      if(_mul_5_source_busy) begin
        _mul_5_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_5_fsm_1 = 1;
  localparam _mul_5_fsm_2 = 2;
  localparam _mul_5_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_fsm <= _mul_5_fsm_init;
      _mul_5_source_start <= 0;
      _mul_5_source_busy <= 0;
      _mul_5_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_5_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_5_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_5_stream_oready && _tmp_417) begin
        _mul_5_stream_ivalid <= 1;
      end 
      if(_mul_5_stream_oready && 1'd0) begin
        _mul_5_stream_ivalid <= 0;
      end 
      case(_mul_5_fsm)
        _mul_5_fsm_init: begin
          if(_mul_5_run_flag) begin
            _mul_5_source_start <= 1;
          end 
          if(_mul_5_run_flag) begin
            _mul_5_fsm <= _mul_5_fsm_1;
          end 
        end
        _mul_5_fsm_1: begin
          if(_mul_5_source_start && _mul_5_stream_oready) begin
            _mul_5_source_start <= 0;
            _mul_5_source_busy <= 1;
          end 
          if(_mul_5_source_start && _mul_5_stream_oready) begin
            _mul_5_fsm <= _mul_5_fsm_2;
          end 
        end
        _mul_5_fsm_2: begin
          if(_mul_5_stream_oready) begin
            _mul_5_fsm <= _mul_5_fsm_3;
          end 
        end
        _mul_5_fsm_3: begin
          if(_mul_5_stream_oready && 1'd0) begin
            _mul_5_source_busy <= 0;
          end 
          if(_mul_5_stream_oready && 1'd0 && _mul_5_run_flag) begin
            _mul_5_source_start <= 1;
          end 
          if(_mul_5_stream_oready && 1'd0) begin
            _mul_5_fsm <= _mul_5_fsm_init;
          end 
          if(_mul_5_stream_oready && 1'd0 && _mul_5_run_flag) begin
            _mul_5_fsm <= _mul_5_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_x_source_ram_renable <= 0;
      _mul_6_x_source_fifo_deq <= 0;
      _mul_6_x_idle <= 1;
      _mul_6_y_source_ram_renable <= 0;
      _mul_6_y_source_fifo_deq <= 0;
      _mul_6_y_idle <= 1;
      _mul_6_rshift_source_ram_renable <= 0;
      _mul_6_rshift_source_fifo_deq <= 0;
      _mul_6_rshift_idle <= 1;
      _mul_6_z_sink_wenable <= 0;
      _mul_6_z_sink_fifo_enq <= 0;
      __mul_6_stream_ivalid_1 <= 0;
      __mul_6_stream_ivalid_2 <= 0;
      __mul_6_stream_ivalid_3 <= 0;
      __mul_6_stream_ivalid_4 <= 0;
      __mul_6_stream_ivalid_5 <= 0;
      __mul_6_stream_ivalid_6 <= 0;
      __mul_6_stream_ivalid_7 <= 0;
      __mul_6_stream_ivalid_8 <= 0;
      _greaterthan_data_136 <= 0;
      _minus_data_138 <= 0;
      _greatereq_data_149 <= 0;
      __delay_data_698__variable_133 <= 0;
      __delay_data_701__variable_134 <= 0;
      __delay_data_704__variable_135 <= 0;
      _sll_data_140 <= 0;
      __delay_data_695_greaterthan_136 <= 0;
      __delay_data_696_greatereq_149 <= 0;
      __delay_data_699__delay_698__variable_133 <= 0;
      __delay_data_702__delay_701__variable_134 <= 0;
      __delay_data_705__delay_704__variable_135 <= 0;
      _cond_data_146 <= 0;
      __delay_data_697__delay_696_greatereq_149 <= 0;
      __delay_data_700__delay_699__delay_698__variable_133 <= 0;
      __delay_data_703__delay_702__delay_701__variable_134 <= 0;
      __delay_data_706__delay_705__delay_704__variable_135 <= 0;
      __muladd_madd_odata_reg_152 <= 0;
      __delay_data_707__delay_706__delay_705____variable_135 <= 0;
      __delay_data_708__delay_707__delay_706____variable_135 <= 0;
      __delay_data_709__delay_708__delay_707____variable_135 <= 0;
      __delay_data_710__delay_709__delay_708____variable_135 <= 0;
      _sra_data_153 <= 0;
      __variable_wdata_133 <= 0;
      __variable_wdata_134 <= 0;
      __variable_wdata_135 <= 0;
      _tmp_449 <= 0;
      _tmp_450 <= 0;
      _tmp_451 <= 0;
      _tmp_452 <= 0;
      _tmp_453 <= 0;
      _tmp_454 <= 0;
      _tmp_455 <= 0;
      _tmp_456 <= 0;
      _tmp_457 <= 0;
      _tmp_458 <= 0;
      _tmp_459 <= 0;
      _tmp_460 <= 0;
      _tmp_461 <= 0;
      _tmp_462 <= 0;
      _tmp_463 <= 0;
      _tmp_464 <= 0;
      _tmp_465 <= 0;
      _tmp_466 <= 0;
      _tmp_467 <= 0;
      _tmp_468 <= 0;
      _tmp_469 <= 0;
      _tmp_470 <= 0;
      _tmp_471 <= 0;
      _tmp_472 <= 0;
      _tmp_473 <= 0;
      _tmp_474 <= 0;
      _tmp_475 <= 0;
      _tmp_476 <= 0;
      _tmp_477 <= 0;
      _tmp_478 <= 0;
      _tmp_479 <= 0;
      _tmp_480 <= 0;
      _tmp_481 <= 0;
      _tmp_482 <= 0;
      _mul_6_busy_reg <= 0;
    end else begin
      if(_mul_6_stream_oready) begin
        _mul_6_x_source_ram_renable <= 0;
        _mul_6_x_source_fifo_deq <= 0;
      end 
      _mul_6_x_idle <= _mul_6_x_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_y_source_ram_renable <= 0;
        _mul_6_y_source_fifo_deq <= 0;
      end 
      _mul_6_y_idle <= _mul_6_y_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_rshift_source_ram_renable <= 0;
        _mul_6_rshift_source_fifo_deq <= 0;
      end 
      _mul_6_rshift_idle <= _mul_6_rshift_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_z_sink_wenable <= 0;
        _mul_6_z_sink_fifo_enq <= 0;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_1 <= _mul_6_stream_ivalid;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_2 <= __mul_6_stream_ivalid_1;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_3 <= __mul_6_stream_ivalid_2;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_4 <= __mul_6_stream_ivalid_3;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_5 <= __mul_6_stream_ivalid_4;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_6 <= __mul_6_stream_ivalid_5;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_7 <= __mul_6_stream_ivalid_6;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_8 <= __mul_6_stream_ivalid_7;
      end 
      if(_mul_6_stream_oready) begin
        _greaterthan_data_136 <= mul_6_rshift_data > 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        _minus_data_138 <= mul_6_rshift_data - 2'sd1;
      end 
      if(_mul_6_stream_oready) begin
        _greatereq_data_149 <= mul_6_x_data >= 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_698__variable_133 <= mul_6_x_data;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_701__variable_134 <= mul_6_y_data;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_704__variable_135 <= mul_6_rshift_data;
      end 
      if(_mul_6_stream_oready) begin
        _sll_data_140 <= 2'sd1 << _minus_data_138;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_695_greaterthan_136 <= _greaterthan_data_136;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_696_greatereq_149 <= _greatereq_data_149;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_699__delay_698__variable_133 <= __delay_data_698__variable_133;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_702__delay_701__variable_134 <= __delay_data_701__variable_134;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_705__delay_704__variable_135 <= __delay_data_704__variable_135;
      end 
      if(_mul_6_stream_oready) begin
        _cond_data_146 <= (__delay_data_695_greaterthan_136)? _sll_data_140 : 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_697__delay_696_greatereq_149 <= __delay_data_696_greatereq_149;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_700__delay_699__delay_698__variable_133 <= __delay_data_699__delay_698__variable_133;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_703__delay_702__delay_701__variable_134 <= __delay_data_702__delay_701__variable_134;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_706__delay_705__delay_704__variable_135 <= __delay_data_705__delay_704__variable_135;
      end 
      if(_mul_6_stream_oready) begin
        __muladd_madd_odata_reg_152 <= __muladd_madd_odata_152;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_707__delay_706__delay_705____variable_135 <= __delay_data_706__delay_705__delay_704__variable_135;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_708__delay_707__delay_706____variable_135 <= __delay_data_707__delay_706__delay_705____variable_135;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_709__delay_708__delay_707____variable_135 <= __delay_data_708__delay_707__delay_706____variable_135;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_710__delay_709__delay_708____variable_135 <= __delay_data_709__delay_708__delay_707____variable_135;
      end 
      if(_mul_6_stream_oready) begin
        _sra_data_153 <= __muladd_data_152 >>> __delay_data_710__delay_709__delay_708____variable_135;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_133 <= _cond_data_626;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_134 <= __delay_data_882_reinterpretcast_595;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_135 <= _plus_data_711;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_449 <= _mul_6_source_start;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_450 <= _tmp_449;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_451 <= _tmp_450;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_452 <= _mul_6_source_start;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_453 <= _tmp_452;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_454 <= _tmp_453;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_455 <= _tmp_454;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_456 <= _tmp_455;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_457 <= _tmp_456;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_458 <= _tmp_457;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_459 <= _tmp_458;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_460 <= _tmp_459;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_461 <= _tmp_460;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_462 <= _mul_6_source_stop;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_463 <= _tmp_462;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_464 <= _tmp_463;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_465 <= _tmp_464;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_466 <= _tmp_465;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_467 <= _tmp_466;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_468 <= _tmp_467;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_469 <= _tmp_468;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_470 <= _tmp_469;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_471 <= _tmp_470;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_472 <= _mul_6_source_busy;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_473 <= _tmp_472;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_474 <= _tmp_473;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_475 <= _tmp_474;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_476 <= _tmp_475;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_477 <= _tmp_476;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_478 <= _tmp_477;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_479 <= _tmp_478;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_480 <= _tmp_479;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_481 <= _tmp_480;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_482 <= _mul_6_sink_busy;
      end 
      if(!_mul_6_sink_busy && _tmp_482) begin
        _mul_6_busy_reg <= 0;
      end 
      if(_mul_6_source_busy) begin
        _mul_6_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_6_fsm_1 = 1;
  localparam _mul_6_fsm_2 = 2;
  localparam _mul_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_fsm <= _mul_6_fsm_init;
      _mul_6_source_start <= 0;
      _mul_6_source_busy <= 0;
      _mul_6_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_6_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_6_stream_oready && _tmp_451) begin
        _mul_6_stream_ivalid <= 1;
      end 
      if(_mul_6_stream_oready && 1'd0) begin
        _mul_6_stream_ivalid <= 0;
      end 
      case(_mul_6_fsm)
        _mul_6_fsm_init: begin
          if(_mul_6_run_flag) begin
            _mul_6_source_start <= 1;
          end 
          if(_mul_6_run_flag) begin
            _mul_6_fsm <= _mul_6_fsm_1;
          end 
        end
        _mul_6_fsm_1: begin
          if(_mul_6_source_start && _mul_6_stream_oready) begin
            _mul_6_source_start <= 0;
            _mul_6_source_busy <= 1;
          end 
          if(_mul_6_source_start && _mul_6_stream_oready) begin
            _mul_6_fsm <= _mul_6_fsm_2;
          end 
        end
        _mul_6_fsm_2: begin
          if(_mul_6_stream_oready) begin
            _mul_6_fsm <= _mul_6_fsm_3;
          end 
        end
        _mul_6_fsm_3: begin
          if(_mul_6_stream_oready && 1'd0) begin
            _mul_6_source_busy <= 0;
          end 
          if(_mul_6_stream_oready && 1'd0 && _mul_6_run_flag) begin
            _mul_6_source_start <= 1;
          end 
          if(_mul_6_stream_oready && 1'd0) begin
            _mul_6_fsm <= _mul_6_fsm_init;
          end 
          if(_mul_6_stream_oready && 1'd0 && _mul_6_run_flag) begin
            _mul_6_fsm <= _mul_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_x_source_ram_renable <= 0;
      _mul_7_x_source_fifo_deq <= 0;
      _mul_7_x_idle <= 1;
      _mul_7_y_source_ram_renable <= 0;
      _mul_7_y_source_fifo_deq <= 0;
      _mul_7_y_idle <= 1;
      _mul_7_rshift_source_ram_renable <= 0;
      _mul_7_rshift_source_fifo_deq <= 0;
      _mul_7_rshift_idle <= 1;
      _mul_7_z_sink_wenable <= 0;
      _mul_7_z_sink_fifo_enq <= 0;
      __mul_7_stream_ivalid_1 <= 0;
      __mul_7_stream_ivalid_2 <= 0;
      __mul_7_stream_ivalid_3 <= 0;
      __mul_7_stream_ivalid_4 <= 0;
      __mul_7_stream_ivalid_5 <= 0;
      __mul_7_stream_ivalid_6 <= 0;
      __mul_7_stream_ivalid_7 <= 0;
      __mul_7_stream_ivalid_8 <= 0;
      _greaterthan_data_157 <= 0;
      _minus_data_159 <= 0;
      _greatereq_data_170 <= 0;
      __delay_data_717__variable_154 <= 0;
      __delay_data_720__variable_155 <= 0;
      __delay_data_723__variable_156 <= 0;
      _sll_data_161 <= 0;
      __delay_data_714_greaterthan_157 <= 0;
      __delay_data_715_greatereq_170 <= 0;
      __delay_data_718__delay_717__variable_154 <= 0;
      __delay_data_721__delay_720__variable_155 <= 0;
      __delay_data_724__delay_723__variable_156 <= 0;
      _cond_data_167 <= 0;
      __delay_data_716__delay_715_greatereq_170 <= 0;
      __delay_data_719__delay_718__delay_717__variable_154 <= 0;
      __delay_data_722__delay_721__delay_720__variable_155 <= 0;
      __delay_data_725__delay_724__delay_723__variable_156 <= 0;
      __muladd_madd_odata_reg_173 <= 0;
      __delay_data_726__delay_725__delay_724____variable_156 <= 0;
      __delay_data_727__delay_726__delay_725____variable_156 <= 0;
      __delay_data_728__delay_727__delay_726____variable_156 <= 0;
      __delay_data_729__delay_728__delay_727____variable_156 <= 0;
      _sra_data_174 <= 0;
      __variable_wdata_154 <= 0;
      __variable_wdata_155 <= 0;
      __variable_wdata_156 <= 0;
      _tmp_483 <= 0;
      _tmp_484 <= 0;
      _tmp_485 <= 0;
      _tmp_486 <= 0;
      _tmp_487 <= 0;
      _tmp_488 <= 0;
      _tmp_489 <= 0;
      _tmp_490 <= 0;
      _tmp_491 <= 0;
      _tmp_492 <= 0;
      _tmp_493 <= 0;
      _tmp_494 <= 0;
      _tmp_495 <= 0;
      _tmp_496 <= 0;
      _tmp_497 <= 0;
      _tmp_498 <= 0;
      _tmp_499 <= 0;
      _tmp_500 <= 0;
      _tmp_501 <= 0;
      _tmp_502 <= 0;
      _tmp_503 <= 0;
      _tmp_504 <= 0;
      _tmp_505 <= 0;
      _tmp_506 <= 0;
      _tmp_507 <= 0;
      _tmp_508 <= 0;
      _tmp_509 <= 0;
      _tmp_510 <= 0;
      _tmp_511 <= 0;
      _tmp_512 <= 0;
      _tmp_513 <= 0;
      _tmp_514 <= 0;
      _tmp_515 <= 0;
      _tmp_516 <= 0;
      _mul_7_busy_reg <= 0;
    end else begin
      if(_mul_7_stream_oready) begin
        _mul_7_x_source_ram_renable <= 0;
        _mul_7_x_source_fifo_deq <= 0;
      end 
      _mul_7_x_idle <= _mul_7_x_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_y_source_ram_renable <= 0;
        _mul_7_y_source_fifo_deq <= 0;
      end 
      _mul_7_y_idle <= _mul_7_y_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_rshift_source_ram_renable <= 0;
        _mul_7_rshift_source_fifo_deq <= 0;
      end 
      _mul_7_rshift_idle <= _mul_7_rshift_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_z_sink_wenable <= 0;
        _mul_7_z_sink_fifo_enq <= 0;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_1 <= _mul_7_stream_ivalid;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_2 <= __mul_7_stream_ivalid_1;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_3 <= __mul_7_stream_ivalid_2;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_4 <= __mul_7_stream_ivalid_3;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_5 <= __mul_7_stream_ivalid_4;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_6 <= __mul_7_stream_ivalid_5;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_7 <= __mul_7_stream_ivalid_6;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_8 <= __mul_7_stream_ivalid_7;
      end 
      if(_mul_7_stream_oready) begin
        _greaterthan_data_157 <= mul_7_rshift_data > 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        _minus_data_159 <= mul_7_rshift_data - 2'sd1;
      end 
      if(_mul_7_stream_oready) begin
        _greatereq_data_170 <= mul_7_x_data >= 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_717__variable_154 <= mul_7_x_data;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_720__variable_155 <= mul_7_y_data;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_723__variable_156 <= mul_7_rshift_data;
      end 
      if(_mul_7_stream_oready) begin
        _sll_data_161 <= 2'sd1 << _minus_data_159;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_714_greaterthan_157 <= _greaterthan_data_157;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_715_greatereq_170 <= _greatereq_data_170;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_718__delay_717__variable_154 <= __delay_data_717__variable_154;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_721__delay_720__variable_155 <= __delay_data_720__variable_155;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_724__delay_723__variable_156 <= __delay_data_723__variable_156;
      end 
      if(_mul_7_stream_oready) begin
        _cond_data_167 <= (__delay_data_714_greaterthan_157)? _sll_data_161 : 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_716__delay_715_greatereq_170 <= __delay_data_715_greatereq_170;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_719__delay_718__delay_717__variable_154 <= __delay_data_718__delay_717__variable_154;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_722__delay_721__delay_720__variable_155 <= __delay_data_721__delay_720__variable_155;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_725__delay_724__delay_723__variable_156 <= __delay_data_724__delay_723__variable_156;
      end 
      if(_mul_7_stream_oready) begin
        __muladd_madd_odata_reg_173 <= __muladd_madd_odata_173;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_726__delay_725__delay_724____variable_156 <= __delay_data_725__delay_724__delay_723__variable_156;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_727__delay_726__delay_725____variable_156 <= __delay_data_726__delay_725__delay_724____variable_156;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_728__delay_727__delay_726____variable_156 <= __delay_data_727__delay_726__delay_725____variable_156;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_729__delay_728__delay_727____variable_156 <= __delay_data_728__delay_727__delay_726____variable_156;
      end 
      if(_mul_7_stream_oready) begin
        _sra_data_174 <= __muladd_data_173 >>> __delay_data_729__delay_728__delay_727____variable_156;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_154 <= _cond_data_628;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_155 <= __delay_data_884_reinterpretcast_596;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_156 <= _plus_data_730;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_483 <= _mul_7_source_start;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_484 <= _tmp_483;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_485 <= _tmp_484;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_486 <= _mul_7_source_start;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_487 <= _tmp_486;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_488 <= _tmp_487;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_489 <= _tmp_488;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_490 <= _tmp_489;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_491 <= _tmp_490;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_492 <= _tmp_491;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_493 <= _tmp_492;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_494 <= _tmp_493;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_495 <= _tmp_494;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_496 <= _mul_7_source_stop;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_497 <= _tmp_496;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_498 <= _tmp_497;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_499 <= _tmp_498;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_500 <= _tmp_499;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_501 <= _tmp_500;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_502 <= _tmp_501;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_503 <= _tmp_502;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_504 <= _tmp_503;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_505 <= _tmp_504;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_506 <= _mul_7_source_busy;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_507 <= _tmp_506;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_508 <= _tmp_507;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_509 <= _tmp_508;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_510 <= _tmp_509;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_511 <= _tmp_510;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_512 <= _tmp_511;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_513 <= _tmp_512;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_514 <= _tmp_513;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_515 <= _tmp_514;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_516 <= _mul_7_sink_busy;
      end 
      if(!_mul_7_sink_busy && _tmp_516) begin
        _mul_7_busy_reg <= 0;
      end 
      if(_mul_7_source_busy) begin
        _mul_7_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_7_fsm_1 = 1;
  localparam _mul_7_fsm_2 = 2;
  localparam _mul_7_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_fsm <= _mul_7_fsm_init;
      _mul_7_source_start <= 0;
      _mul_7_source_busy <= 0;
      _mul_7_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_7_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_7_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_7_stream_oready && _tmp_485) begin
        _mul_7_stream_ivalid <= 1;
      end 
      if(_mul_7_stream_oready && 1'd0) begin
        _mul_7_stream_ivalid <= 0;
      end 
      case(_mul_7_fsm)
        _mul_7_fsm_init: begin
          if(_mul_7_run_flag) begin
            _mul_7_source_start <= 1;
          end 
          if(_mul_7_run_flag) begin
            _mul_7_fsm <= _mul_7_fsm_1;
          end 
        end
        _mul_7_fsm_1: begin
          if(_mul_7_source_start && _mul_7_stream_oready) begin
            _mul_7_source_start <= 0;
            _mul_7_source_busy <= 1;
          end 
          if(_mul_7_source_start && _mul_7_stream_oready) begin
            _mul_7_fsm <= _mul_7_fsm_2;
          end 
        end
        _mul_7_fsm_2: begin
          if(_mul_7_stream_oready) begin
            _mul_7_fsm <= _mul_7_fsm_3;
          end 
        end
        _mul_7_fsm_3: begin
          if(_mul_7_stream_oready && 1'd0) begin
            _mul_7_source_busy <= 0;
          end 
          if(_mul_7_stream_oready && 1'd0 && _mul_7_run_flag) begin
            _mul_7_source_start <= 1;
          end 
          if(_mul_7_stream_oready && 1'd0) begin
            _mul_7_fsm <= _mul_7_fsm_init;
          end 
          if(_mul_7_stream_oready && 1'd0 && _mul_7_run_flag) begin
            _mul_7_fsm <= _mul_7_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_x_source_ram_renable <= 0;
      _mul_8_x_source_fifo_deq <= 0;
      _mul_8_x_idle <= 1;
      _mul_8_y_source_ram_renable <= 0;
      _mul_8_y_source_fifo_deq <= 0;
      _mul_8_y_idle <= 1;
      _mul_8_rshift_source_ram_renable <= 0;
      _mul_8_rshift_source_fifo_deq <= 0;
      _mul_8_rshift_idle <= 1;
      _mul_8_z_sink_wenable <= 0;
      _mul_8_z_sink_fifo_enq <= 0;
      __mul_8_stream_ivalid_1 <= 0;
      __mul_8_stream_ivalid_2 <= 0;
      __mul_8_stream_ivalid_3 <= 0;
      __mul_8_stream_ivalid_4 <= 0;
      __mul_8_stream_ivalid_5 <= 0;
      __mul_8_stream_ivalid_6 <= 0;
      __mul_8_stream_ivalid_7 <= 0;
      __mul_8_stream_ivalid_8 <= 0;
      _greaterthan_data_178 <= 0;
      _minus_data_180 <= 0;
      _greatereq_data_191 <= 0;
      __delay_data_736__variable_175 <= 0;
      __delay_data_739__variable_176 <= 0;
      __delay_data_742__variable_177 <= 0;
      _sll_data_182 <= 0;
      __delay_data_733_greaterthan_178 <= 0;
      __delay_data_734_greatereq_191 <= 0;
      __delay_data_737__delay_736__variable_175 <= 0;
      __delay_data_740__delay_739__variable_176 <= 0;
      __delay_data_743__delay_742__variable_177 <= 0;
      _cond_data_188 <= 0;
      __delay_data_735__delay_734_greatereq_191 <= 0;
      __delay_data_738__delay_737__delay_736__variable_175 <= 0;
      __delay_data_741__delay_740__delay_739__variable_176 <= 0;
      __delay_data_744__delay_743__delay_742__variable_177 <= 0;
      __muladd_madd_odata_reg_194 <= 0;
      __delay_data_745__delay_744__delay_743____variable_177 <= 0;
      __delay_data_746__delay_745__delay_744____variable_177 <= 0;
      __delay_data_747__delay_746__delay_745____variable_177 <= 0;
      __delay_data_748__delay_747__delay_746____variable_177 <= 0;
      _sra_data_195 <= 0;
      __variable_wdata_175 <= 0;
      __variable_wdata_176 <= 0;
      __variable_wdata_177 <= 0;
      _tmp_517 <= 0;
      _tmp_518 <= 0;
      _tmp_519 <= 0;
      _tmp_520 <= 0;
      _tmp_521 <= 0;
      _tmp_522 <= 0;
      _tmp_523 <= 0;
      _tmp_524 <= 0;
      _tmp_525 <= 0;
      _tmp_526 <= 0;
      _tmp_527 <= 0;
      _tmp_528 <= 0;
      _tmp_529 <= 0;
      _tmp_530 <= 0;
      _tmp_531 <= 0;
      _tmp_532 <= 0;
      _tmp_533 <= 0;
      _tmp_534 <= 0;
      _tmp_535 <= 0;
      _tmp_536 <= 0;
      _tmp_537 <= 0;
      _tmp_538 <= 0;
      _tmp_539 <= 0;
      _tmp_540 <= 0;
      _tmp_541 <= 0;
      _tmp_542 <= 0;
      _tmp_543 <= 0;
      _tmp_544 <= 0;
      _tmp_545 <= 0;
      _tmp_546 <= 0;
      _tmp_547 <= 0;
      _tmp_548 <= 0;
      _tmp_549 <= 0;
      _tmp_550 <= 0;
      _mul_8_busy_reg <= 0;
    end else begin
      if(_mul_8_stream_oready) begin
        _mul_8_x_source_ram_renable <= 0;
        _mul_8_x_source_fifo_deq <= 0;
      end 
      _mul_8_x_idle <= _mul_8_x_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_y_source_ram_renable <= 0;
        _mul_8_y_source_fifo_deq <= 0;
      end 
      _mul_8_y_idle <= _mul_8_y_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_rshift_source_ram_renable <= 0;
        _mul_8_rshift_source_fifo_deq <= 0;
      end 
      _mul_8_rshift_idle <= _mul_8_rshift_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_z_sink_wenable <= 0;
        _mul_8_z_sink_fifo_enq <= 0;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_1 <= _mul_8_stream_ivalid;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_2 <= __mul_8_stream_ivalid_1;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_3 <= __mul_8_stream_ivalid_2;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_4 <= __mul_8_stream_ivalid_3;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_5 <= __mul_8_stream_ivalid_4;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_6 <= __mul_8_stream_ivalid_5;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_7 <= __mul_8_stream_ivalid_6;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_8 <= __mul_8_stream_ivalid_7;
      end 
      if(_mul_8_stream_oready) begin
        _greaterthan_data_178 <= mul_8_rshift_data > 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        _minus_data_180 <= mul_8_rshift_data - 2'sd1;
      end 
      if(_mul_8_stream_oready) begin
        _greatereq_data_191 <= mul_8_x_data >= 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_736__variable_175 <= mul_8_x_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_739__variable_176 <= mul_8_y_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_742__variable_177 <= mul_8_rshift_data;
      end 
      if(_mul_8_stream_oready) begin
        _sll_data_182 <= 2'sd1 << _minus_data_180;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_733_greaterthan_178 <= _greaterthan_data_178;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_734_greatereq_191 <= _greatereq_data_191;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_737__delay_736__variable_175 <= __delay_data_736__variable_175;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_740__delay_739__variable_176 <= __delay_data_739__variable_176;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_743__delay_742__variable_177 <= __delay_data_742__variable_177;
      end 
      if(_mul_8_stream_oready) begin
        _cond_data_188 <= (__delay_data_733_greaterthan_178)? _sll_data_182 : 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_735__delay_734_greatereq_191 <= __delay_data_734_greatereq_191;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_738__delay_737__delay_736__variable_175 <= __delay_data_737__delay_736__variable_175;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_741__delay_740__delay_739__variable_176 <= __delay_data_740__delay_739__variable_176;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_744__delay_743__delay_742__variable_177 <= __delay_data_743__delay_742__variable_177;
      end 
      if(_mul_8_stream_oready) begin
        __muladd_madd_odata_reg_194 <= __muladd_madd_odata_194;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_745__delay_744__delay_743____variable_177 <= __delay_data_744__delay_743__delay_742__variable_177;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_746__delay_745__delay_744____variable_177 <= __delay_data_745__delay_744__delay_743____variable_177;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_747__delay_746__delay_745____variable_177 <= __delay_data_746__delay_745__delay_744____variable_177;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_748__delay_747__delay_746____variable_177 <= __delay_data_747__delay_746__delay_745____variable_177;
      end 
      if(_mul_8_stream_oready) begin
        _sra_data_195 <= __muladd_data_194 >>> __delay_data_748__delay_747__delay_746____variable_177;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_175 <= _cond_data_630;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_176 <= __delay_data_886_reinterpretcast_597;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_177 <= _plus_data_749;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_517 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_518 <= _tmp_517;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_519 <= _tmp_518;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_520 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_521 <= _tmp_520;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_522 <= _tmp_521;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_523 <= _tmp_522;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_524 <= _tmp_523;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_525 <= _tmp_524;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_526 <= _tmp_525;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_527 <= _tmp_526;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_528 <= _tmp_527;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_529 <= _tmp_528;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_530 <= _mul_8_source_stop;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_531 <= _tmp_530;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_532 <= _tmp_531;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_533 <= _tmp_532;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_534 <= _tmp_533;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_535 <= _tmp_534;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_536 <= _tmp_535;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_537 <= _tmp_536;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_538 <= _tmp_537;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_539 <= _tmp_538;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_540 <= _mul_8_source_busy;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_541 <= _tmp_540;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_542 <= _tmp_541;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_543 <= _tmp_542;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_544 <= _tmp_543;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_545 <= _tmp_544;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_546 <= _tmp_545;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_547 <= _tmp_546;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_548 <= _tmp_547;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_549 <= _tmp_548;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_550 <= _mul_8_sink_busy;
      end 
      if(!_mul_8_sink_busy && _tmp_550) begin
        _mul_8_busy_reg <= 0;
      end 
      if(_mul_8_source_busy) begin
        _mul_8_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_8_fsm_1 = 1;
  localparam _mul_8_fsm_2 = 2;
  localparam _mul_8_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_fsm <= _mul_8_fsm_init;
      _mul_8_source_start <= 0;
      _mul_8_source_busy <= 0;
      _mul_8_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_8_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_8_stream_oready && _tmp_519) begin
        _mul_8_stream_ivalid <= 1;
      end 
      if(_mul_8_stream_oready && 1'd0) begin
        _mul_8_stream_ivalid <= 0;
      end 
      case(_mul_8_fsm)
        _mul_8_fsm_init: begin
          if(_mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
        _mul_8_fsm_1: begin
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_source_start <= 0;
            _mul_8_source_busy <= 1;
          end 
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_2;
          end 
        end
        _mul_8_fsm_2: begin
          if(_mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_3;
          end 
        end
        _mul_8_fsm_3: begin
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_source_busy <= 0;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_fsm <= _mul_8_fsm_init;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_x_source_ram_renable <= 0;
      _mul_9_x_source_fifo_deq <= 0;
      _mul_9_x_idle <= 1;
      _mul_9_y_source_ram_renable <= 0;
      _mul_9_y_source_fifo_deq <= 0;
      _mul_9_y_idle <= 1;
      _mul_9_rshift_source_ram_renable <= 0;
      _mul_9_rshift_source_fifo_deq <= 0;
      _mul_9_rshift_idle <= 1;
      _mul_9_z_sink_wenable <= 0;
      _mul_9_z_sink_fifo_enq <= 0;
      __mul_9_stream_ivalid_1 <= 0;
      __mul_9_stream_ivalid_2 <= 0;
      __mul_9_stream_ivalid_3 <= 0;
      __mul_9_stream_ivalid_4 <= 0;
      __mul_9_stream_ivalid_5 <= 0;
      __mul_9_stream_ivalid_6 <= 0;
      __mul_9_stream_ivalid_7 <= 0;
      __mul_9_stream_ivalid_8 <= 0;
      _greaterthan_data_199 <= 0;
      _minus_data_201 <= 0;
      _greatereq_data_212 <= 0;
      __delay_data_755__variable_196 <= 0;
      __delay_data_758__variable_197 <= 0;
      __delay_data_761__variable_198 <= 0;
      _sll_data_203 <= 0;
      __delay_data_752_greaterthan_199 <= 0;
      __delay_data_753_greatereq_212 <= 0;
      __delay_data_756__delay_755__variable_196 <= 0;
      __delay_data_759__delay_758__variable_197 <= 0;
      __delay_data_762__delay_761__variable_198 <= 0;
      _cond_data_209 <= 0;
      __delay_data_754__delay_753_greatereq_212 <= 0;
      __delay_data_757__delay_756__delay_755__variable_196 <= 0;
      __delay_data_760__delay_759__delay_758__variable_197 <= 0;
      __delay_data_763__delay_762__delay_761__variable_198 <= 0;
      __muladd_madd_odata_reg_215 <= 0;
      __delay_data_764__delay_763__delay_762____variable_198 <= 0;
      __delay_data_765__delay_764__delay_763____variable_198 <= 0;
      __delay_data_766__delay_765__delay_764____variable_198 <= 0;
      __delay_data_767__delay_766__delay_765____variable_198 <= 0;
      _sra_data_216 <= 0;
      __variable_wdata_196 <= 0;
      __variable_wdata_197 <= 0;
      __variable_wdata_198 <= 0;
      _tmp_551 <= 0;
      _tmp_552 <= 0;
      _tmp_553 <= 0;
      _tmp_554 <= 0;
      _tmp_555 <= 0;
      _tmp_556 <= 0;
      _tmp_557 <= 0;
      _tmp_558 <= 0;
      _tmp_559 <= 0;
      _tmp_560 <= 0;
      _tmp_561 <= 0;
      _tmp_562 <= 0;
      _tmp_563 <= 0;
      _tmp_564 <= 0;
      _tmp_565 <= 0;
      _tmp_566 <= 0;
      _tmp_567 <= 0;
      _tmp_568 <= 0;
      _tmp_569 <= 0;
      _tmp_570 <= 0;
      _tmp_571 <= 0;
      _tmp_572 <= 0;
      _tmp_573 <= 0;
      _tmp_574 <= 0;
      _tmp_575 <= 0;
      _tmp_576 <= 0;
      _tmp_577 <= 0;
      _tmp_578 <= 0;
      _tmp_579 <= 0;
      _tmp_580 <= 0;
      _tmp_581 <= 0;
      _tmp_582 <= 0;
      _tmp_583 <= 0;
      _tmp_584 <= 0;
      _mul_9_busy_reg <= 0;
    end else begin
      if(_mul_9_stream_oready) begin
        _mul_9_x_source_ram_renable <= 0;
        _mul_9_x_source_fifo_deq <= 0;
      end 
      _mul_9_x_idle <= _mul_9_x_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_y_source_ram_renable <= 0;
        _mul_9_y_source_fifo_deq <= 0;
      end 
      _mul_9_y_idle <= _mul_9_y_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_rshift_source_ram_renable <= 0;
        _mul_9_rshift_source_fifo_deq <= 0;
      end 
      _mul_9_rshift_idle <= _mul_9_rshift_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_z_sink_wenable <= 0;
        _mul_9_z_sink_fifo_enq <= 0;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_1 <= _mul_9_stream_ivalid;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_2 <= __mul_9_stream_ivalid_1;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_3 <= __mul_9_stream_ivalid_2;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_4 <= __mul_9_stream_ivalid_3;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_5 <= __mul_9_stream_ivalid_4;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_6 <= __mul_9_stream_ivalid_5;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_7 <= __mul_9_stream_ivalid_6;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_8 <= __mul_9_stream_ivalid_7;
      end 
      if(_mul_9_stream_oready) begin
        _greaterthan_data_199 <= mul_9_rshift_data > 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        _minus_data_201 <= mul_9_rshift_data - 2'sd1;
      end 
      if(_mul_9_stream_oready) begin
        _greatereq_data_212 <= mul_9_x_data >= 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_755__variable_196 <= mul_9_x_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_758__variable_197 <= mul_9_y_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_761__variable_198 <= mul_9_rshift_data;
      end 
      if(_mul_9_stream_oready) begin
        _sll_data_203 <= 2'sd1 << _minus_data_201;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_752_greaterthan_199 <= _greaterthan_data_199;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_753_greatereq_212 <= _greatereq_data_212;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_756__delay_755__variable_196 <= __delay_data_755__variable_196;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_759__delay_758__variable_197 <= __delay_data_758__variable_197;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_762__delay_761__variable_198 <= __delay_data_761__variable_198;
      end 
      if(_mul_9_stream_oready) begin
        _cond_data_209 <= (__delay_data_752_greaterthan_199)? _sll_data_203 : 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_754__delay_753_greatereq_212 <= __delay_data_753_greatereq_212;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_757__delay_756__delay_755__variable_196 <= __delay_data_756__delay_755__variable_196;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_760__delay_759__delay_758__variable_197 <= __delay_data_759__delay_758__variable_197;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_763__delay_762__delay_761__variable_198 <= __delay_data_762__delay_761__variable_198;
      end 
      if(_mul_9_stream_oready) begin
        __muladd_madd_odata_reg_215 <= __muladd_madd_odata_215;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_764__delay_763__delay_762____variable_198 <= __delay_data_763__delay_762__delay_761__variable_198;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_765__delay_764__delay_763____variable_198 <= __delay_data_764__delay_763__delay_762____variable_198;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_766__delay_765__delay_764____variable_198 <= __delay_data_765__delay_764__delay_763____variable_198;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_767__delay_766__delay_765____variable_198 <= __delay_data_766__delay_765__delay_764____variable_198;
      end 
      if(_mul_9_stream_oready) begin
        _sra_data_216 <= __muladd_data_215 >>> __delay_data_767__delay_766__delay_765____variable_198;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_196 <= _cond_data_632;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_197 <= __delay_data_888_reinterpretcast_598;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_198 <= _plus_data_768;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_551 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_552 <= _tmp_551;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_553 <= _tmp_552;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_554 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_555 <= _tmp_554;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_556 <= _tmp_555;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_557 <= _tmp_556;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_558 <= _tmp_557;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_559 <= _tmp_558;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_560 <= _tmp_559;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_561 <= _tmp_560;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_562 <= _tmp_561;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_563 <= _tmp_562;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_564 <= _mul_9_source_stop;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_565 <= _tmp_564;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_566 <= _tmp_565;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_567 <= _tmp_566;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_568 <= _tmp_567;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_569 <= _tmp_568;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_570 <= _tmp_569;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_571 <= _tmp_570;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_572 <= _tmp_571;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_573 <= _tmp_572;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_574 <= _mul_9_source_busy;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_575 <= _tmp_574;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_576 <= _tmp_575;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_577 <= _tmp_576;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_578 <= _tmp_577;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_579 <= _tmp_578;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_580 <= _tmp_579;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_581 <= _tmp_580;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_582 <= _tmp_581;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_583 <= _tmp_582;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_584 <= _mul_9_sink_busy;
      end 
      if(!_mul_9_sink_busy && _tmp_584) begin
        _mul_9_busy_reg <= 0;
      end 
      if(_mul_9_source_busy) begin
        _mul_9_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_9_fsm_1 = 1;
  localparam _mul_9_fsm_2 = 2;
  localparam _mul_9_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_fsm <= _mul_9_fsm_init;
      _mul_9_source_start <= 0;
      _mul_9_source_busy <= 0;
      _mul_9_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_9_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_9_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_9_stream_oready && _tmp_553) begin
        _mul_9_stream_ivalid <= 1;
      end 
      if(_mul_9_stream_oready && 1'd0) begin
        _mul_9_stream_ivalid <= 0;
      end 
      case(_mul_9_fsm)
        _mul_9_fsm_init: begin
          if(_mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
        _mul_9_fsm_1: begin
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_source_start <= 0;
            _mul_9_source_busy <= 1;
          end 
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_2;
          end 
        end
        _mul_9_fsm_2: begin
          if(_mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_3;
          end 
        end
        _mul_9_fsm_3: begin
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_source_busy <= 0;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_fsm <= _mul_9_fsm_init;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_x_source_ram_renable <= 0;
      _mul_10_x_source_fifo_deq <= 0;
      _mul_10_x_idle <= 1;
      _mul_10_y_source_ram_renable <= 0;
      _mul_10_y_source_fifo_deq <= 0;
      _mul_10_y_idle <= 1;
      _mul_10_rshift_source_ram_renable <= 0;
      _mul_10_rshift_source_fifo_deq <= 0;
      _mul_10_rshift_idle <= 1;
      _mul_10_z_sink_wenable <= 0;
      _mul_10_z_sink_fifo_enq <= 0;
      __mul_10_stream_ivalid_1 <= 0;
      __mul_10_stream_ivalid_2 <= 0;
      __mul_10_stream_ivalid_3 <= 0;
      __mul_10_stream_ivalid_4 <= 0;
      __mul_10_stream_ivalid_5 <= 0;
      __mul_10_stream_ivalid_6 <= 0;
      __mul_10_stream_ivalid_7 <= 0;
      __mul_10_stream_ivalid_8 <= 0;
      _greaterthan_data_220 <= 0;
      _minus_data_222 <= 0;
      _greatereq_data_233 <= 0;
      __delay_data_774__variable_217 <= 0;
      __delay_data_777__variable_218 <= 0;
      __delay_data_780__variable_219 <= 0;
      _sll_data_224 <= 0;
      __delay_data_771_greaterthan_220 <= 0;
      __delay_data_772_greatereq_233 <= 0;
      __delay_data_775__delay_774__variable_217 <= 0;
      __delay_data_778__delay_777__variable_218 <= 0;
      __delay_data_781__delay_780__variable_219 <= 0;
      _cond_data_230 <= 0;
      __delay_data_773__delay_772_greatereq_233 <= 0;
      __delay_data_776__delay_775__delay_774__variable_217 <= 0;
      __delay_data_779__delay_778__delay_777__variable_218 <= 0;
      __delay_data_782__delay_781__delay_780__variable_219 <= 0;
      __muladd_madd_odata_reg_236 <= 0;
      __delay_data_783__delay_782__delay_781____variable_219 <= 0;
      __delay_data_784__delay_783__delay_782____variable_219 <= 0;
      __delay_data_785__delay_784__delay_783____variable_219 <= 0;
      __delay_data_786__delay_785__delay_784____variable_219 <= 0;
      _sra_data_237 <= 0;
      __variable_wdata_217 <= 0;
      __variable_wdata_218 <= 0;
      __variable_wdata_219 <= 0;
      _tmp_585 <= 0;
      _tmp_586 <= 0;
      _tmp_587 <= 0;
      _tmp_588 <= 0;
      _tmp_589 <= 0;
      _tmp_590 <= 0;
      _tmp_591 <= 0;
      _tmp_592 <= 0;
      _tmp_593 <= 0;
      _tmp_594 <= 0;
      _tmp_595 <= 0;
      _tmp_596 <= 0;
      _tmp_597 <= 0;
      _tmp_598 <= 0;
      _tmp_599 <= 0;
      _tmp_600 <= 0;
      _tmp_601 <= 0;
      _tmp_602 <= 0;
      _tmp_603 <= 0;
      _tmp_604 <= 0;
      _tmp_605 <= 0;
      _tmp_606 <= 0;
      _tmp_607 <= 0;
      _tmp_608 <= 0;
      _tmp_609 <= 0;
      _tmp_610 <= 0;
      _tmp_611 <= 0;
      _tmp_612 <= 0;
      _tmp_613 <= 0;
      _tmp_614 <= 0;
      _tmp_615 <= 0;
      _tmp_616 <= 0;
      _tmp_617 <= 0;
      _tmp_618 <= 0;
      _mul_10_busy_reg <= 0;
    end else begin
      if(_mul_10_stream_oready) begin
        _mul_10_x_source_ram_renable <= 0;
        _mul_10_x_source_fifo_deq <= 0;
      end 
      _mul_10_x_idle <= _mul_10_x_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_y_source_ram_renable <= 0;
        _mul_10_y_source_fifo_deq <= 0;
      end 
      _mul_10_y_idle <= _mul_10_y_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_rshift_source_ram_renable <= 0;
        _mul_10_rshift_source_fifo_deq <= 0;
      end 
      _mul_10_rshift_idle <= _mul_10_rshift_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_z_sink_wenable <= 0;
        _mul_10_z_sink_fifo_enq <= 0;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_1 <= _mul_10_stream_ivalid;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_2 <= __mul_10_stream_ivalid_1;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_3 <= __mul_10_stream_ivalid_2;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_4 <= __mul_10_stream_ivalid_3;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_5 <= __mul_10_stream_ivalid_4;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_6 <= __mul_10_stream_ivalid_5;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_7 <= __mul_10_stream_ivalid_6;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_8 <= __mul_10_stream_ivalid_7;
      end 
      if(_mul_10_stream_oready) begin
        _greaterthan_data_220 <= mul_10_rshift_data > 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        _minus_data_222 <= mul_10_rshift_data - 2'sd1;
      end 
      if(_mul_10_stream_oready) begin
        _greatereq_data_233 <= mul_10_x_data >= 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_774__variable_217 <= mul_10_x_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_777__variable_218 <= mul_10_y_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_780__variable_219 <= mul_10_rshift_data;
      end 
      if(_mul_10_stream_oready) begin
        _sll_data_224 <= 2'sd1 << _minus_data_222;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_771_greaterthan_220 <= _greaterthan_data_220;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_772_greatereq_233 <= _greatereq_data_233;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_775__delay_774__variable_217 <= __delay_data_774__variable_217;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_778__delay_777__variable_218 <= __delay_data_777__variable_218;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_781__delay_780__variable_219 <= __delay_data_780__variable_219;
      end 
      if(_mul_10_stream_oready) begin
        _cond_data_230 <= (__delay_data_771_greaterthan_220)? _sll_data_224 : 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_773__delay_772_greatereq_233 <= __delay_data_772_greatereq_233;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_776__delay_775__delay_774__variable_217 <= __delay_data_775__delay_774__variable_217;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_779__delay_778__delay_777__variable_218 <= __delay_data_778__delay_777__variable_218;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_782__delay_781__delay_780__variable_219 <= __delay_data_781__delay_780__variable_219;
      end 
      if(_mul_10_stream_oready) begin
        __muladd_madd_odata_reg_236 <= __muladd_madd_odata_236;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_783__delay_782__delay_781____variable_219 <= __delay_data_782__delay_781__delay_780__variable_219;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_784__delay_783__delay_782____variable_219 <= __delay_data_783__delay_782__delay_781____variable_219;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_785__delay_784__delay_783____variable_219 <= __delay_data_784__delay_783__delay_782____variable_219;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_786__delay_785__delay_784____variable_219 <= __delay_data_785__delay_784__delay_783____variable_219;
      end 
      if(_mul_10_stream_oready) begin
        _sra_data_237 <= __muladd_data_236 >>> __delay_data_786__delay_785__delay_784____variable_219;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_217 <= _cond_data_634;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_218 <= __delay_data_890_reinterpretcast_599;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_219 <= _plus_data_787;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_585 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_586 <= _tmp_585;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_587 <= _tmp_586;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_588 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_589 <= _tmp_588;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_590 <= _tmp_589;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_591 <= _tmp_590;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_592 <= _tmp_591;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_593 <= _tmp_592;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_594 <= _tmp_593;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_595 <= _tmp_594;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_596 <= _tmp_595;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_597 <= _tmp_596;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_598 <= _mul_10_source_stop;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_599 <= _tmp_598;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_600 <= _tmp_599;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_601 <= _tmp_600;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_602 <= _tmp_601;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_603 <= _tmp_602;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_604 <= _tmp_603;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_605 <= _tmp_604;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_606 <= _tmp_605;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_607 <= _tmp_606;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_608 <= _mul_10_source_busy;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_609 <= _tmp_608;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_610 <= _tmp_609;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_611 <= _tmp_610;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_612 <= _tmp_611;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_613 <= _tmp_612;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_614 <= _tmp_613;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_615 <= _tmp_614;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_616 <= _tmp_615;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_617 <= _tmp_616;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_618 <= _mul_10_sink_busy;
      end 
      if(!_mul_10_sink_busy && _tmp_618) begin
        _mul_10_busy_reg <= 0;
      end 
      if(_mul_10_source_busy) begin
        _mul_10_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_10_fsm_1 = 1;
  localparam _mul_10_fsm_2 = 2;
  localparam _mul_10_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_fsm <= _mul_10_fsm_init;
      _mul_10_source_start <= 0;
      _mul_10_source_busy <= 0;
      _mul_10_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_10_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_10_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_10_stream_oready && _tmp_587) begin
        _mul_10_stream_ivalid <= 1;
      end 
      if(_mul_10_stream_oready && 1'd0) begin
        _mul_10_stream_ivalid <= 0;
      end 
      case(_mul_10_fsm)
        _mul_10_fsm_init: begin
          if(_mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
        _mul_10_fsm_1: begin
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_source_start <= 0;
            _mul_10_source_busy <= 1;
          end 
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_2;
          end 
        end
        _mul_10_fsm_2: begin
          if(_mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_3;
          end 
        end
        _mul_10_fsm_3: begin
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_source_busy <= 0;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_fsm <= _mul_10_fsm_init;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_x_source_ram_renable <= 0;
      _mul_11_x_source_fifo_deq <= 0;
      _mul_11_x_idle <= 1;
      _mul_11_y_source_ram_renable <= 0;
      _mul_11_y_source_fifo_deq <= 0;
      _mul_11_y_idle <= 1;
      _mul_11_rshift_source_ram_renable <= 0;
      _mul_11_rshift_source_fifo_deq <= 0;
      _mul_11_rshift_idle <= 1;
      _mul_11_z_sink_wenable <= 0;
      _mul_11_z_sink_fifo_enq <= 0;
      __mul_11_stream_ivalid_1 <= 0;
      __mul_11_stream_ivalid_2 <= 0;
      __mul_11_stream_ivalid_3 <= 0;
      __mul_11_stream_ivalid_4 <= 0;
      __mul_11_stream_ivalid_5 <= 0;
      __mul_11_stream_ivalid_6 <= 0;
      __mul_11_stream_ivalid_7 <= 0;
      __mul_11_stream_ivalid_8 <= 0;
      _greaterthan_data_241 <= 0;
      _minus_data_243 <= 0;
      _greatereq_data_254 <= 0;
      __delay_data_793__variable_238 <= 0;
      __delay_data_796__variable_239 <= 0;
      __delay_data_799__variable_240 <= 0;
      _sll_data_245 <= 0;
      __delay_data_790_greaterthan_241 <= 0;
      __delay_data_791_greatereq_254 <= 0;
      __delay_data_794__delay_793__variable_238 <= 0;
      __delay_data_797__delay_796__variable_239 <= 0;
      __delay_data_800__delay_799__variable_240 <= 0;
      _cond_data_251 <= 0;
      __delay_data_792__delay_791_greatereq_254 <= 0;
      __delay_data_795__delay_794__delay_793__variable_238 <= 0;
      __delay_data_798__delay_797__delay_796__variable_239 <= 0;
      __delay_data_801__delay_800__delay_799__variable_240 <= 0;
      __muladd_madd_odata_reg_257 <= 0;
      __delay_data_802__delay_801__delay_800____variable_240 <= 0;
      __delay_data_803__delay_802__delay_801____variable_240 <= 0;
      __delay_data_804__delay_803__delay_802____variable_240 <= 0;
      __delay_data_805__delay_804__delay_803____variable_240 <= 0;
      _sra_data_258 <= 0;
      __variable_wdata_238 <= 0;
      __variable_wdata_239 <= 0;
      __variable_wdata_240 <= 0;
      _tmp_619 <= 0;
      _tmp_620 <= 0;
      _tmp_621 <= 0;
      _tmp_622 <= 0;
      _tmp_623 <= 0;
      _tmp_624 <= 0;
      _tmp_625 <= 0;
      _tmp_626 <= 0;
      _tmp_627 <= 0;
      _tmp_628 <= 0;
      _tmp_629 <= 0;
      _tmp_630 <= 0;
      _tmp_631 <= 0;
      _tmp_632 <= 0;
      _tmp_633 <= 0;
      _tmp_634 <= 0;
      _tmp_635 <= 0;
      _tmp_636 <= 0;
      _tmp_637 <= 0;
      _tmp_638 <= 0;
      _tmp_639 <= 0;
      _tmp_640 <= 0;
      _tmp_641 <= 0;
      _tmp_642 <= 0;
      _tmp_643 <= 0;
      _tmp_644 <= 0;
      _tmp_645 <= 0;
      _tmp_646 <= 0;
      _tmp_647 <= 0;
      _tmp_648 <= 0;
      _tmp_649 <= 0;
      _tmp_650 <= 0;
      _tmp_651 <= 0;
      _tmp_652 <= 0;
      _mul_11_busy_reg <= 0;
    end else begin
      if(_mul_11_stream_oready) begin
        _mul_11_x_source_ram_renable <= 0;
        _mul_11_x_source_fifo_deq <= 0;
      end 
      _mul_11_x_idle <= _mul_11_x_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_y_source_ram_renable <= 0;
        _mul_11_y_source_fifo_deq <= 0;
      end 
      _mul_11_y_idle <= _mul_11_y_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_rshift_source_ram_renable <= 0;
        _mul_11_rshift_source_fifo_deq <= 0;
      end 
      _mul_11_rshift_idle <= _mul_11_rshift_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_z_sink_wenable <= 0;
        _mul_11_z_sink_fifo_enq <= 0;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_1 <= _mul_11_stream_ivalid;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_2 <= __mul_11_stream_ivalid_1;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_3 <= __mul_11_stream_ivalid_2;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_4 <= __mul_11_stream_ivalid_3;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_5 <= __mul_11_stream_ivalid_4;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_6 <= __mul_11_stream_ivalid_5;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_7 <= __mul_11_stream_ivalid_6;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_8 <= __mul_11_stream_ivalid_7;
      end 
      if(_mul_11_stream_oready) begin
        _greaterthan_data_241 <= mul_11_rshift_data > 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        _minus_data_243 <= mul_11_rshift_data - 2'sd1;
      end 
      if(_mul_11_stream_oready) begin
        _greatereq_data_254 <= mul_11_x_data >= 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_793__variable_238 <= mul_11_x_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_796__variable_239 <= mul_11_y_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_799__variable_240 <= mul_11_rshift_data;
      end 
      if(_mul_11_stream_oready) begin
        _sll_data_245 <= 2'sd1 << _minus_data_243;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_790_greaterthan_241 <= _greaterthan_data_241;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_791_greatereq_254 <= _greatereq_data_254;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_794__delay_793__variable_238 <= __delay_data_793__variable_238;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_797__delay_796__variable_239 <= __delay_data_796__variable_239;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_800__delay_799__variable_240 <= __delay_data_799__variable_240;
      end 
      if(_mul_11_stream_oready) begin
        _cond_data_251 <= (__delay_data_790_greaterthan_241)? _sll_data_245 : 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_792__delay_791_greatereq_254 <= __delay_data_791_greatereq_254;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_795__delay_794__delay_793__variable_238 <= __delay_data_794__delay_793__variable_238;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_798__delay_797__delay_796__variable_239 <= __delay_data_797__delay_796__variable_239;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_801__delay_800__delay_799__variable_240 <= __delay_data_800__delay_799__variable_240;
      end 
      if(_mul_11_stream_oready) begin
        __muladd_madd_odata_reg_257 <= __muladd_madd_odata_257;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_802__delay_801__delay_800____variable_240 <= __delay_data_801__delay_800__delay_799__variable_240;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_803__delay_802__delay_801____variable_240 <= __delay_data_802__delay_801__delay_800____variable_240;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_804__delay_803__delay_802____variable_240 <= __delay_data_803__delay_802__delay_801____variable_240;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_805__delay_804__delay_803____variable_240 <= __delay_data_804__delay_803__delay_802____variable_240;
      end 
      if(_mul_11_stream_oready) begin
        _sra_data_258 <= __muladd_data_257 >>> __delay_data_805__delay_804__delay_803____variable_240;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_238 <= _cond_data_636;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_239 <= __delay_data_892_reinterpretcast_600;
      end 
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        __variable_wdata_240 <= _plus_data_806;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_619 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_620 <= _tmp_619;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_621 <= _tmp_620;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_622 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_623 <= _tmp_622;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_624 <= _tmp_623;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_625 <= _tmp_624;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_626 <= _tmp_625;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_627 <= _tmp_626;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_628 <= _tmp_627;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_629 <= _tmp_628;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_630 <= _tmp_629;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_631 <= _tmp_630;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_632 <= _mul_11_source_stop;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_633 <= _tmp_632;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_634 <= _tmp_633;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_635 <= _tmp_634;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_636 <= _tmp_635;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_637 <= _tmp_636;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_638 <= _tmp_637;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_639 <= _tmp_638;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_640 <= _tmp_639;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_641 <= _tmp_640;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_642 <= _mul_11_source_busy;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_643 <= _tmp_642;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_644 <= _tmp_643;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_645 <= _tmp_644;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_646 <= _tmp_645;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_647 <= _tmp_646;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_648 <= _tmp_647;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_649 <= _tmp_648;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_650 <= _tmp_649;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_651 <= _tmp_650;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_652 <= _mul_11_sink_busy;
      end 
      if(!_mul_11_sink_busy && _tmp_652) begin
        _mul_11_busy_reg <= 0;
      end 
      if(_mul_11_source_busy) begin
        _mul_11_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_11_fsm_1 = 1;
  localparam _mul_11_fsm_2 = 2;
  localparam _mul_11_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_fsm <= _mul_11_fsm_init;
      _mul_11_source_start <= 0;
      _mul_11_source_busy <= 0;
      _mul_11_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_2_stream_ivalid_1 && _stream_conv2d_2_stream_oready) begin
        _mul_11_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_busy) begin
        _mul_11_source_busy <= _stream_conv2d_2_source_busy;
      end 
      if(_mul_11_stream_oready && _tmp_621) begin
        _mul_11_stream_ivalid <= 1;
      end 
      if(_mul_11_stream_oready && 1'd0) begin
        _mul_11_stream_ivalid <= 0;
      end 
      case(_mul_11_fsm)
        _mul_11_fsm_init: begin
          if(_mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
        _mul_11_fsm_1: begin
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_source_start <= 0;
            _mul_11_source_busy <= 1;
          end 
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_2;
          end 
        end
        _mul_11_fsm_2: begin
          if(_mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_3;
          end 
        end
        _mul_11_fsm_3: begin
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_source_busy <= 0;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_fsm <= _mul_11_fsm_init;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_7_source_ram_renable <= 0;
      _stream_conv2d_2_source_7_source_fifo_deq <= 0;
      _stream_conv2d_2_source_7_idle <= 1;
      _stream_conv2d_2_source_9_source_ram_renable <= 0;
      _stream_conv2d_2_source_9_source_fifo_deq <= 0;
      _stream_conv2d_2_source_9_idle <= 1;
      _stream_conv2d_2_source_11_source_ram_renable <= 0;
      _stream_conv2d_2_source_11_source_fifo_deq <= 0;
      _stream_conv2d_2_source_11_idle <= 1;
      _stream_conv2d_2_source_13_source_ram_renable <= 0;
      _stream_conv2d_2_source_13_source_fifo_deq <= 0;
      _stream_conv2d_2_source_13_idle <= 1;
      _stream_conv2d_2_source_15_source_ram_renable <= 0;
      _stream_conv2d_2_source_15_source_fifo_deq <= 0;
      _stream_conv2d_2_source_15_idle <= 1;
      _stream_conv2d_2_source_20_source_ram_renable <= 0;
      _stream_conv2d_2_source_20_source_fifo_deq <= 0;
      _stream_conv2d_2_source_20_idle <= 1;
      _stream_conv2d_2_source_21_source_ram_renable <= 0;
      _stream_conv2d_2_source_21_source_fifo_deq <= 0;
      _stream_conv2d_2_source_21_idle <= 1;
      _stream_conv2d_2_source_22_source_ram_renable <= 0;
      _stream_conv2d_2_source_22_source_fifo_deq <= 0;
      _stream_conv2d_2_source_22_idle <= 1;
      _stream_conv2d_2_source_23_source_ram_renable <= 0;
      _stream_conv2d_2_source_23_source_fifo_deq <= 0;
      _stream_conv2d_2_source_23_idle <= 1;
      _stream_conv2d_2_source_24_source_ram_renable <= 0;
      _stream_conv2d_2_source_24_source_fifo_deq <= 0;
      _stream_conv2d_2_source_24_idle <= 1;
      _stream_conv2d_2_source_25_source_ram_renable <= 0;
      _stream_conv2d_2_source_25_source_fifo_deq <= 0;
      _stream_conv2d_2_source_25_idle <= 1;
      _stream_conv2d_2_source_26_source_ram_renable <= 0;
      _stream_conv2d_2_source_26_source_fifo_deq <= 0;
      _stream_conv2d_2_source_26_idle <= 1;
      _stream_conv2d_2_source_27_source_ram_renable <= 0;
      _stream_conv2d_2_source_27_source_fifo_deq <= 0;
      _stream_conv2d_2_source_27_idle <= 1;
      _stream_conv2d_2_source_28_source_ram_renable <= 0;
      _stream_conv2d_2_source_28_source_fifo_deq <= 0;
      _stream_conv2d_2_source_28_idle <= 1;
      _stream_conv2d_2_source_29_source_ram_renable <= 0;
      _stream_conv2d_2_source_29_source_fifo_deq <= 0;
      _stream_conv2d_2_source_29_idle <= 1;
      _stream_conv2d_2_source_30_source_ram_renable <= 0;
      _stream_conv2d_2_source_30_source_fifo_deq <= 0;
      _stream_conv2d_2_source_30_idle <= 1;
      _stream_conv2d_2_source_31_source_ram_renable <= 0;
      _stream_conv2d_2_source_31_source_fifo_deq <= 0;
      _stream_conv2d_2_source_31_idle <= 1;
      _stream_conv2d_2_source_32_source_ram_renable <= 0;
      _stream_conv2d_2_source_32_source_fifo_deq <= 0;
      _stream_conv2d_2_source_32_idle <= 1;
      _stream_conv2d_2_source_33_source_ram_renable <= 0;
      _stream_conv2d_2_source_33_source_fifo_deq <= 0;
      _stream_conv2d_2_source_33_idle <= 1;
      _stream_conv2d_2_source_34_source_ram_renable <= 0;
      _stream_conv2d_2_source_34_source_fifo_deq <= 0;
      _stream_conv2d_2_source_34_idle <= 1;
      _stream_conv2d_2_source_35_source_ram_renable <= 0;
      _stream_conv2d_2_source_35_source_fifo_deq <= 0;
      _stream_conv2d_2_source_35_idle <= 1;
      _stream_conv2d_2_source_36_source_ram_renable <= 0;
      _stream_conv2d_2_source_36_source_fifo_deq <= 0;
      _stream_conv2d_2_source_36_idle <= 1;
      _stream_conv2d_2_source_37_source_ram_renable <= 0;
      _stream_conv2d_2_source_37_source_fifo_deq <= 0;
      _stream_conv2d_2_source_37_idle <= 1;
      _stream_conv2d_2_sink_50_sink_wenable <= 0;
      _stream_conv2d_2_sink_50_sink_fifo_enq <= 0;
      _stream_conv2d_2_sink_51_sink_wenable <= 0;
      _stream_conv2d_2_sink_51_sink_fifo_enq <= 0;
      __stream_conv2d_2_stream_ivalid_1 <= 0;
      __stream_conv2d_2_stream_ivalid_2 <= 0;
      __stream_conv2d_2_stream_ivalid_3 <= 0;
      __stream_conv2d_2_stream_ivalid_4 <= 0;
      __stream_conv2d_2_stream_ivalid_5 <= 0;
      __stream_conv2d_2_stream_ivalid_6 <= 0;
      __stream_conv2d_2_stream_ivalid_7 <= 0;
      __stream_conv2d_2_stream_ivalid_8 <= 0;
      __stream_conv2d_2_stream_ivalid_9 <= 0;
      __stream_conv2d_2_stream_ivalid_10 <= 0;
      __stream_conv2d_2_stream_ivalid_11 <= 0;
      __stream_conv2d_2_stream_ivalid_12 <= 0;
      __stream_conv2d_2_stream_ivalid_13 <= 0;
      __stream_conv2d_2_stream_ivalid_14 <= 0;
      __stream_conv2d_2_stream_ivalid_15 <= 0;
      __stream_conv2d_2_stream_ivalid_16 <= 0;
      __stream_conv2d_2_stream_ivalid_17 <= 0;
      __stream_conv2d_2_stream_ivalid_18 <= 0;
      __stream_conv2d_2_stream_ivalid_19 <= 0;
      __stream_conv2d_2_stream_ivalid_20 <= 0;
      __stream_conv2d_2_stream_ivalid_21 <= 0;
      __stream_conv2d_2_stream_ivalid_22 <= 0;
      __stream_conv2d_2_stream_ivalid_23 <= 0;
      __stream_conv2d_2_stream_ivalid_24 <= 0;
      __stream_conv2d_2_stream_ivalid_25 <= 0;
      __stream_conv2d_2_stream_ivalid_26 <= 0;
      __stream_conv2d_2_stream_ivalid_27 <= 0;
      __stream_conv2d_2_stream_ivalid_28 <= 0;
      __stream_conv2d_2_stream_ivalid_29 <= 0;
      _eq_data_322 <= 0;
      _eq_data_326 <= 0;
      _eq_data_329 <= 0;
      _eq_data_332 <= 0;
      _eq_data_336 <= 0;
      _eq_data_339 <= 0;
      _eq_data_342 <= 0;
      _eq_data_346 <= 0;
      _eq_data_349 <= 0;
      _eq_data_352 <= 0;
      _eq_data_356 <= 0;
      _eq_data_359 <= 0;
      _eq_data_362 <= 0;
      _eq_data_366 <= 0;
      _eq_data_369 <= 0;
      _eq_data_372 <= 0;
      _eq_data_376 <= 0;
      _eq_data_379 <= 0;
      _eq_data_382 <= 0;
      _eq_data_386 <= 0;
      _eq_data_389 <= 0;
      _eq_data_392 <= 0;
      _eq_data_396 <= 0;
      _eq_data_399 <= 0;
      _eq_data_402 <= 0;
      _eq_data_406 <= 0;
      _eq_data_409 <= 0;
      _eq_data_412 <= 0;
      _eq_data_416 <= 0;
      _eq_data_419 <= 0;
      _eq_data_422 <= 0;
      _eq_data_426 <= 0;
      _eq_data_429 <= 0;
      _eq_data_432 <= 0;
      _eq_data_436 <= 0;
      _eq_data_439 <= 0;
      _eq_data_442 <= 0;
      _eq_data_446 <= 0;
      _eq_data_449 <= 0;
      _eq_data_452 <= 0;
      _eq_data_456 <= 0;
      _eq_data_459 <= 0;
      _eq_data_462 <= 0;
      _eq_data_466 <= 0;
      _eq_data_469 <= 0;
      _eq_data_472 <= 0;
      _eq_data_476 <= 0;
      _eq_data_479 <= 0;
      _eq_data_482 <= 0;
      _eq_data_486 <= 0;
      _eq_data_489 <= 0;
      _eq_data_492 <= 0;
      _eq_data_496 <= 0;
      _eq_data_499 <= 0;
      _plus_data_654 <= 0;
      _plus_data_673 <= 0;
      _plus_data_692 <= 0;
      _plus_data_711 <= 0;
      _plus_data_730 <= 0;
      _plus_data_749 <= 0;
      _plus_data_768 <= 0;
      _plus_data_787 <= 0;
      _plus_data_806 <= 0;
      _plus_data_822 <= 0;
      _plus_data_841 <= 0;
      __delay_data_866__variable_315 <= 0;
      __delay_data_867__variable_314 <= 0;
      __delay_data_868__variable_313 <= 0;
      __delay_data_869__variable_318 <= 0;
      __delay_data_870__variable_317 <= 0;
      __delay_data_871__variable_316 <= 0;
      __delay_data_872__variable_321 <= 0;
      __delay_data_873__variable_320 <= 0;
      __delay_data_874__variable_319 <= 0;
      __delay_data_875_pointer_601 <= 0;
      __delay_data_876_reinterpretcast_592 <= 0;
      __delay_data_877_pointer_603 <= 0;
      __delay_data_878_reinterpretcast_593 <= 0;
      __delay_data_879_pointer_605 <= 0;
      __delay_data_880_reinterpretcast_594 <= 0;
      __delay_data_881_pointer_607 <= 0;
      __delay_data_882_reinterpretcast_595 <= 0;
      __delay_data_883_pointer_609 <= 0;
      __delay_data_884_reinterpretcast_596 <= 0;
      __delay_data_885_pointer_611 <= 0;
      __delay_data_886_reinterpretcast_597 <= 0;
      __delay_data_887_pointer_613 <= 0;
      __delay_data_888_reinterpretcast_598 <= 0;
      __delay_data_889_pointer_615 <= 0;
      __delay_data_890_reinterpretcast_599 <= 0;
      __delay_data_891_pointer_617 <= 0;
      __delay_data_892_reinterpretcast_600 <= 0;
      __delay_data_893__variable_264 <= 0;
      __delay_data_918__variable_259 <= 0;
      __delay_data_931_cond_280 <= 0;
      __delay_data_950_cond_287 <= 0;
      __delay_data_894__delay_893__variable_264 <= 0;
      __delay_data_906_plus_822 <= 0;
      __delay_data_919__delay_918__variable_259 <= 0;
      __delay_data_932__delay_931_cond_280 <= 0;
      __delay_data_951__delay_950_cond_287 <= 0;
      __delay_data_970_plus_841 <= 0;
      __delay_data_895__delay_894__delay_893__variable_264 <= 0;
      __delay_data_907__delay_906_plus_822 <= 0;
      __delay_data_920__delay_919__delay_918__variable_259 <= 0;
      __delay_data_933__delay_932__delay_931_cond_280 <= 0;
      __delay_data_952__delay_951__delay_950_cond_287 <= 0;
      __delay_data_971__delay_970_plus_841 <= 0;
      __delay_data_896__delay_895__delay_894____variable_264 <= 0;
      __delay_data_908__delay_907__delay_906_plus_822 <= 0;
      __delay_data_921__delay_920__delay_919____variable_259 <= 0;
      __delay_data_934__delay_933__delay_932__delay_931_cond_280 <= 0;
      __delay_data_953__delay_952__delay_951__delay_950_cond_287 <= 0;
      __delay_data_972__delay_971__delay_970_plus_841 <= 0;
      __delay_data_897__delay_896__delay_895____variable_264 <= 0;
      __delay_data_909__delay_908__delay_907__delay_906_plus_822 <= 0;
      __delay_data_922__delay_921__delay_920____variable_259 <= 0;
      __delay_data_935__delay_934__delay_933__delay_932___cond_280 <= 0;
      __delay_data_954__delay_953__delay_952__delay_951___cond_287 <= 0;
      __delay_data_973__delay_972__delay_971__delay_970_plus_841 <= 0;
      __delay_data_898__delay_897__delay_896____variable_264 <= 0;
      __delay_data_910__delay_909__delay_908__delay_907___plus_822 <= 0;
      __delay_data_923__delay_922__delay_921____variable_259 <= 0;
      __delay_data_936__delay_935__delay_934__delay_933___cond_280 <= 0;
      __delay_data_955__delay_954__delay_953__delay_952___cond_287 <= 0;
      __delay_data_974__delay_973__delay_972__delay_971___plus_841 <= 0;
      __delay_data_899__delay_898__delay_897____variable_264 <= 0;
      __delay_data_911__delay_910__delay_909__delay_908___plus_822 <= 0;
      __delay_data_924__delay_923__delay_922____variable_259 <= 0;
      __delay_data_937__delay_936__delay_935__delay_934___cond_280 <= 0;
      __delay_data_956__delay_955__delay_954__delay_953___cond_287 <= 0;
      __delay_data_975__delay_974__delay_973__delay_972___plus_841 <= 0;
      __delay_data_900__delay_899__delay_898____variable_264 <= 0;
      __delay_data_912__delay_911__delay_910__delay_909___plus_822 <= 0;
      __delay_data_925__delay_924__delay_923____variable_259 <= 0;
      __delay_data_938__delay_937__delay_936__delay_935___cond_280 <= 0;
      __delay_data_957__delay_956__delay_955__delay_954___cond_287 <= 0;
      __delay_data_976__delay_975__delay_974__delay_973___plus_841 <= 0;
      __delay_data_901__delay_900__delay_899____variable_264 <= 0;
      __delay_data_913__delay_912__delay_911__delay_910___plus_822 <= 0;
      __delay_data_926__delay_925__delay_924____variable_259 <= 0;
      __delay_data_939__delay_938__delay_937__delay_936___cond_280 <= 0;
      __delay_data_958__delay_957__delay_956__delay_955___cond_287 <= 0;
      __delay_data_977__delay_976__delay_975__delay_974___plus_841 <= 0;
      __delay_data_902__delay_901__delay_900____variable_264 <= 0;
      __delay_data_914__delay_913__delay_912__delay_911___plus_822 <= 0;
      __delay_data_927__delay_926__delay_925____variable_259 <= 0;
      __delay_data_940__delay_939__delay_938__delay_937___cond_280 <= 0;
      __delay_data_959__delay_958__delay_957__delay_956___cond_287 <= 0;
      __delay_data_978__delay_977__delay_976__delay_975___plus_841 <= 0;
      __delay_data_903__delay_902__delay_901____variable_264 <= 0;
      __delay_data_915__delay_914__delay_913__delay_912___plus_822 <= 0;
      __delay_data_928__delay_927__delay_926____variable_259 <= 0;
      __delay_data_941__delay_940__delay_939__delay_938___cond_280 <= 0;
      __delay_data_960__delay_959__delay_958__delay_957___cond_287 <= 0;
      __delay_data_979__delay_978__delay_977__delay_976___plus_841 <= 0;
      __delay_data_904__delay_903__delay_902____variable_264 <= 0;
      __delay_data_916__delay_915__delay_914__delay_913___plus_822 <= 0;
      __delay_data_929__delay_928__delay_927____variable_259 <= 0;
      __delay_data_942__delay_941__delay_940__delay_939___cond_280 <= 0;
      __delay_data_961__delay_960__delay_959__delay_958___cond_287 <= 0;
      __delay_data_980__delay_979__delay_978__delay_977___plus_841 <= 0;
      __delay_data_905__delay_904__delay_903____variable_264 <= 0;
      __delay_data_917__delay_916__delay_915__delay_914___plus_822 <= 0;
      __delay_data_930__delay_929__delay_928____variable_259 <= 0;
      __delay_data_943__delay_942__delay_941__delay_940___cond_280 <= 0;
      __delay_data_962__delay_961__delay_960__delay_959___cond_287 <= 0;
      __delay_data_981__delay_980__delay_979__delay_978___plus_841 <= 0;
      __delay_data_944__delay_943__delay_942__delay_941___cond_280 <= 0;
      __delay_data_963__delay_962__delay_961__delay_960___cond_287 <= 0;
      __delay_data_982__delay_981__delay_980__delay_979___plus_841 <= 0;
      __delay_data_945__delay_944__delay_943__delay_942___cond_280 <= 0;
      __delay_data_964__delay_963__delay_962__delay_961___cond_287 <= 0;
      __delay_data_983__delay_982__delay_981__delay_980___plus_841 <= 0;
      __delay_data_946__delay_945__delay_944__delay_943___cond_280 <= 0;
      __delay_data_965__delay_964__delay_963__delay_962___cond_287 <= 0;
      __delay_data_984__delay_983__delay_982__delay_981___plus_841 <= 0;
      __delay_data_947__delay_946__delay_945__delay_944___cond_280 <= 0;
      __delay_data_966__delay_965__delay_964__delay_963___cond_287 <= 0;
      __delay_data_985__delay_984__delay_983__delay_982___plus_841 <= 0;
      __delay_data_948__delay_947__delay_946__delay_945___cond_280 <= 0;
      __delay_data_967__delay_966__delay_965__delay_964___cond_287 <= 0;
      __delay_data_986__delay_985__delay_984__delay_983___plus_841 <= 0;
      __delay_data_949__delay_948__delay_947__delay_946___cond_280 <= 0;
      __delay_data_968__delay_967__delay_966__delay_965___cond_287 <= 0;
      __delay_data_987__delay_986__delay_985__delay_984___plus_841 <= 0;
      _plus_data_825 <= 0;
      __delay_data_969__delay_968__delay_967__delay_966___cond_287 <= 0;
      __delay_data_988__delay_987__delay_986__delay_985___plus_841 <= 0;
      __delay_data_989__substreamoutput_824 <= 0;
      __delay_data_990__delay_989__substreamoutput_824 <= 0;
      __delay_data_991__delay_990__delay_989__substreamoutput_824 <= 0;
      __delay_data_992__delay_991__delay_990____substreamoutput_824 <= 0;
      __delay_data_993__delay_992__delay_991____substreamoutput_824 <= 0;
      __delay_data_994__delay_993__delay_992____substreamoutput_824 <= 0;
      __delay_data_995__delay_994__delay_993____substreamoutput_824 <= 0;
      __delay_data_996__delay_995__delay_994____substreamoutput_824 <= 0;
      __delay_data_997__delay_996__delay_995____substreamoutput_824 <= 0;
      __delay_data_998__delay_997__delay_996____substreamoutput_824 <= 0;
      _stream_conv2d_2_parameter_0_next_parameter_data <= 0;
      __variable_wdata_259 <= 0;
      _stream_conv2d_2_parameter_1_next_parameter_data <= 0;
      __variable_wdata_260 <= 0;
      _stream_conv2d_2_parameter_2_next_parameter_data <= 0;
      __variable_wdata_261 <= 0;
      _stream_conv2d_2_parameter_3_next_parameter_data <= 0;
      __variable_wdata_262 <= 0;
      _stream_conv2d_2_parameter_4_next_parameter_data <= 0;
      __variable_wdata_263 <= 0;
      _stream_conv2d_2_parameter_6_next_parameter_data <= 0;
      __variable_wdata_274 <= 0;
      _stream_conv2d_2_source_7_source_mode <= 5'b0;
      _stream_conv2d_2_source_7_source_empty_data <= 0;
      __variable_wdata_275 <= 0;
      _stream_conv2d_2_parameter_8_next_parameter_data <= 0;
      __variable_wdata_281 <= 0;
      _stream_conv2d_2_source_9_source_mode <= 5'b0;
      _stream_conv2d_2_source_9_source_empty_data <= 0;
      __variable_wdata_282 <= 0;
      _stream_conv2d_2_parameter_10_next_parameter_data <= 0;
      __variable_wdata_288 <= 0;
      _stream_conv2d_2_source_11_source_mode <= 5'b0;
      _stream_conv2d_2_source_11_source_empty_data <= 0;
      __variable_wdata_289 <= 0;
      _stream_conv2d_2_parameter_12_next_parameter_data <= 0;
      __variable_wdata_295 <= 0;
      _stream_conv2d_2_source_13_source_mode <= 5'b0;
      _stream_conv2d_2_source_13_source_empty_data <= 0;
      __variable_wdata_296 <= 0;
      _stream_conv2d_2_parameter_14_next_parameter_data <= 0;
      __variable_wdata_302 <= 0;
      _stream_conv2d_2_source_15_source_mode <= 5'b0;
      _stream_conv2d_2_source_15_source_empty_data <= 0;
      __variable_wdata_303 <= 0;
      _stream_conv2d_2_parameter_16_next_parameter_data <= 0;
      __variable_wdata_309 <= 0;
      _stream_conv2d_2_parameter_17_next_parameter_data <= 0;
      __variable_wdata_310 <= 0;
      _stream_conv2d_2_parameter_18_next_parameter_data <= 0;
      __variable_wdata_311 <= 0;
      _stream_conv2d_2_parameter_19_next_parameter_data <= 0;
      __variable_wdata_312 <= 0;
      _stream_conv2d_2_source_20_source_mode <= 5'b0;
      _stream_conv2d_2_source_20_source_offset <= 0;
      _source_stream_conv2d_2_source_20_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_20_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_20_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_20_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_3 <= 0;
      _stream_conv2d_2_source_20_source_sel <= 0;
      _stream_conv2d_2_source_20_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_20_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_20_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_20_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_20_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_20_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_20_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_20_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_20_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_20_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_20_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_20_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_20_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_313 <= 0;
      _stream_conv2d_2_source_20_source_ram_raddr <= 0;
      _stream_conv2d_2_source_21_source_mode <= 5'b0;
      _stream_conv2d_2_source_21_source_offset <= 0;
      _source_stream_conv2d_2_source_21_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_21_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_21_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_21_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_3 <= 0;
      _stream_conv2d_2_source_21_source_sel <= 0;
      _stream_conv2d_2_source_21_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_21_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_21_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_21_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_21_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_21_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_21_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_21_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_21_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_21_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_21_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_21_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_21_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_314 <= 0;
      _stream_conv2d_2_source_21_source_ram_raddr <= 0;
      _stream_conv2d_2_source_22_source_mode <= 5'b0;
      _stream_conv2d_2_source_22_source_offset <= 0;
      _source_stream_conv2d_2_source_22_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_22_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_22_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_22_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_3 <= 0;
      _stream_conv2d_2_source_22_source_sel <= 0;
      _stream_conv2d_2_source_22_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_22_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_22_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_22_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_22_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_22_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_22_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_22_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_22_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_22_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_22_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_22_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_22_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_315 <= 0;
      _stream_conv2d_2_source_22_source_ram_raddr <= 0;
      _stream_conv2d_2_source_23_source_mode <= 5'b0;
      _stream_conv2d_2_source_23_source_offset <= 0;
      _source_stream_conv2d_2_source_23_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_23_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_23_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_23_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_3 <= 0;
      _stream_conv2d_2_source_23_source_sel <= 0;
      _stream_conv2d_2_source_23_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_23_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_23_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_23_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_23_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_23_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_23_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_23_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_23_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_23_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_23_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_23_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_23_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_23_pat_stride_buf_3 <= 0;
      __variable_wdata_316 <= 0;
      _stream_conv2d_2_source_23_source_ram_raddr <= 0;
      _stream_conv2d_2_source_24_source_mode <= 5'b0;
      _stream_conv2d_2_source_24_source_offset <= 0;
      _source_stream_conv2d_2_source_24_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_24_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_24_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_24_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_3 <= 0;
      _stream_conv2d_2_source_24_source_sel <= 0;
      _stream_conv2d_2_source_24_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_24_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_24_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_24_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_24_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_24_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_24_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_24_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_24_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_24_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_24_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_24_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_24_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_24_pat_stride_buf_3 <= 0;
      __variable_wdata_317 <= 0;
      _stream_conv2d_2_source_24_source_ram_raddr <= 0;
      _stream_conv2d_2_source_25_source_mode <= 5'b0;
      _stream_conv2d_2_source_25_source_offset <= 0;
      _source_stream_conv2d_2_source_25_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_25_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_25_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_25_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_3 <= 0;
      _stream_conv2d_2_source_25_source_sel <= 0;
      _stream_conv2d_2_source_25_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_25_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_25_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_25_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_25_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_25_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_25_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_25_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_25_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_25_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_25_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_25_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_25_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_25_pat_stride_buf_3 <= 0;
      __variable_wdata_318 <= 0;
      _stream_conv2d_2_source_25_source_ram_raddr <= 0;
      _stream_conv2d_2_source_26_source_mode <= 5'b0;
      _stream_conv2d_2_source_26_source_offset <= 0;
      _source_stream_conv2d_2_source_26_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_26_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_26_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_26_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_3 <= 0;
      _stream_conv2d_2_source_26_source_sel <= 0;
      _stream_conv2d_2_source_26_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_26_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_26_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_26_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_26_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_26_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_26_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_26_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_26_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_26_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_26_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_26_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_26_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_26_pat_stride_buf_3 <= 0;
      __variable_wdata_319 <= 0;
      _stream_conv2d_2_source_26_source_ram_raddr <= 0;
      _stream_conv2d_2_source_27_source_mode <= 5'b0;
      _stream_conv2d_2_source_27_source_offset <= 0;
      _source_stream_conv2d_2_source_27_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_27_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_27_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_27_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_3 <= 0;
      _stream_conv2d_2_source_27_source_sel <= 0;
      _stream_conv2d_2_source_27_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_27_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_27_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_27_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_27_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_27_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_27_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_27_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_27_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_27_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_27_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_27_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_27_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_27_pat_stride_buf_3 <= 0;
      __variable_wdata_320 <= 0;
      _stream_conv2d_2_source_27_source_ram_raddr <= 0;
      _stream_conv2d_2_source_28_source_mode <= 5'b0;
      _stream_conv2d_2_source_28_source_offset <= 0;
      _source_stream_conv2d_2_source_28_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_28_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_28_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_28_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_3 <= 0;
      _stream_conv2d_2_source_28_source_sel <= 0;
      _stream_conv2d_2_source_28_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_28_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_28_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_28_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_28_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_28_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_28_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_28_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_28_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_28_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_28_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_28_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_28_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_28_pat_stride_buf_3 <= 0;
      __variable_wdata_321 <= 0;
      _stream_conv2d_2_source_28_source_ram_raddr <= 0;
      _stream_conv2d_2_source_29_source_mode <= 5'b0;
      _stream_conv2d_2_source_29_source_offset <= 0;
      _source_stream_conv2d_2_source_29_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_29_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_29_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_29_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_3 <= 0;
      _stream_conv2d_2_source_29_source_sel <= 0;
      _stream_conv2d_2_source_29_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_29_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_29_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_29_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_29_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_29_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_29_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_29_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_29_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_29_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_29_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_29_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_29_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_29_pat_stride_buf_3 <= 0;
      __variable_wdata_547 <= 0;
      _stream_conv2d_2_source_29_source_ram_raddr <= 0;
      _stream_conv2d_2_source_30_source_mode <= 5'b0;
      _stream_conv2d_2_source_30_source_offset <= 0;
      _source_stream_conv2d_2_source_30_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_30_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_30_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_30_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_3 <= 0;
      _stream_conv2d_2_source_30_source_sel <= 0;
      _stream_conv2d_2_source_30_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_30_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_30_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_30_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_30_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_30_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_30_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_30_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_30_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_30_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_30_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_30_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_30_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_30_pat_stride_buf_3 <= 0;
      __variable_wdata_548 <= 0;
      _stream_conv2d_2_source_30_source_ram_raddr <= 0;
      _stream_conv2d_2_source_31_source_mode <= 5'b0;
      _stream_conv2d_2_source_31_source_offset <= 0;
      _source_stream_conv2d_2_source_31_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_31_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_31_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_31_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_3 <= 0;
      _stream_conv2d_2_source_31_source_sel <= 0;
      _stream_conv2d_2_source_31_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_31_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_31_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_31_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_31_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_31_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_31_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_31_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_31_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_31_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_31_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_31_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_31_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_31_pat_stride_buf_3 <= 0;
      __variable_wdata_549 <= 0;
      _stream_conv2d_2_source_31_source_ram_raddr <= 0;
      _stream_conv2d_2_source_32_source_mode <= 5'b0;
      _stream_conv2d_2_source_32_source_offset <= 0;
      _source_stream_conv2d_2_source_32_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_32_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_32_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_32_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_3 <= 0;
      _stream_conv2d_2_source_32_source_sel <= 0;
      _stream_conv2d_2_source_32_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_32_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_32_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_32_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_32_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_32_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_32_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_32_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_32_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_32_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_32_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_32_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_32_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_32_pat_stride_buf_3 <= 0;
      __variable_wdata_550 <= 0;
      _stream_conv2d_2_source_32_source_ram_raddr <= 0;
      _stream_conv2d_2_source_33_source_mode <= 5'b0;
      _stream_conv2d_2_source_33_source_offset <= 0;
      _source_stream_conv2d_2_source_33_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_33_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_33_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_33_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_3 <= 0;
      _stream_conv2d_2_source_33_source_sel <= 0;
      _stream_conv2d_2_source_33_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_33_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_33_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_33_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_33_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_33_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_33_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_33_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_33_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_33_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_33_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_33_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_33_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_33_pat_stride_buf_3 <= 0;
      __variable_wdata_551 <= 0;
      _stream_conv2d_2_source_33_source_ram_raddr <= 0;
      _stream_conv2d_2_source_34_source_mode <= 5'b0;
      _stream_conv2d_2_source_34_source_offset <= 0;
      _source_stream_conv2d_2_source_34_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_34_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_34_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_34_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_3 <= 0;
      _stream_conv2d_2_source_34_source_sel <= 0;
      _stream_conv2d_2_source_34_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_34_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_34_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_34_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_34_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_34_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_34_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_34_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_34_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_34_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_34_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_34_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_34_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_34_pat_stride_buf_3 <= 0;
      __variable_wdata_552 <= 0;
      _stream_conv2d_2_source_34_source_ram_raddr <= 0;
      _stream_conv2d_2_source_35_source_mode <= 5'b0;
      _stream_conv2d_2_source_35_source_offset <= 0;
      _source_stream_conv2d_2_source_35_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_35_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_35_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_35_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_3 <= 0;
      _stream_conv2d_2_source_35_source_sel <= 0;
      _stream_conv2d_2_source_35_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_35_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_35_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_35_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_35_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_35_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_35_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_35_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_35_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_35_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_35_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_35_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_35_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_35_pat_stride_buf_3 <= 0;
      __variable_wdata_553 <= 0;
      _stream_conv2d_2_source_35_source_ram_raddr <= 0;
      _stream_conv2d_2_source_36_source_mode <= 5'b0;
      _stream_conv2d_2_source_36_source_offset <= 0;
      _source_stream_conv2d_2_source_36_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_36_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_36_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_36_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_3 <= 0;
      _stream_conv2d_2_source_36_source_sel <= 0;
      _stream_conv2d_2_source_36_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_36_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_36_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_36_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_36_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_36_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_36_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_36_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_36_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_36_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_36_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_36_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_36_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_36_pat_stride_buf_3 <= 0;
      __variable_wdata_554 <= 0;
      _stream_conv2d_2_source_36_source_ram_raddr <= 0;
      _stream_conv2d_2_source_37_source_mode <= 5'b0;
      _stream_conv2d_2_source_37_source_offset <= 0;
      _source_stream_conv2d_2_source_37_pat_size_0 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_0 <= 0;
      _source_stream_conv2d_2_source_37_pat_size_1 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_1 <= 0;
      _source_stream_conv2d_2_source_37_pat_size_2 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_2 <= 0;
      _source_stream_conv2d_2_source_37_pat_size_3 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_3 <= 0;
      _stream_conv2d_2_source_37_source_sel <= 0;
      _stream_conv2d_2_source_37_source_offset_buf <= 0;
      _source_stream_conv2d_2_source_37_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_2_source_37_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_2_source_37_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_2_source_37_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_2_source_37_pat_count_0 <= 0;
      _source_stream_conv2d_2_source_37_pat_count_1 <= 0;
      _source_stream_conv2d_2_source_37_pat_count_2 <= 0;
      _source_stream_conv2d_2_source_37_pat_count_3 <= 0;
      _source_stream_conv2d_2_source_37_pat_size_buf_0 <= 0;
      _source_stream_conv2d_2_source_37_pat_size_buf_1 <= 0;
      _source_stream_conv2d_2_source_37_pat_size_buf_2 <= 0;
      _source_stream_conv2d_2_source_37_pat_size_buf_3 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_2_source_37_pat_stride_buf_3 <= 0;
      __variable_wdata_555 <= 0;
      _stream_conv2d_2_source_37_source_ram_raddr <= 0;
      _tmp_251 <= 0;
      _tmp_252 <= 0;
      _tmp_253 <= 0;
      _tmp_254 <= 0;
      _tmp_255 <= 0;
      _tmp_256 <= 0;
      _tmp_257 <= 0;
      _tmp_258 <= 0;
      _tmp_259 <= 0;
      _tmp_260 <= 0;
      _tmp_261 <= 0;
      _tmp_262 <= 0;
      _tmp_263 <= 0;
      _tmp_264 <= 0;
      _tmp_265 <= 0;
      _tmp_266 <= 0;
      _tmp_267 <= 0;
      _tmp_268 <= 0;
      _tmp_269 <= 0;
      _tmp_270 <= 0;
      _tmp_271 <= 0;
      _tmp_272 <= 0;
      _tmp_273 <= 0;
      _tmp_274 <= 0;
      _tmp_275 <= 0;
      _tmp_276 <= 0;
      _tmp_277 <= 0;
      _tmp_278 <= 0;
      _tmp_279 <= 0;
      _tmp_280 <= 0;
      _tmp_281 <= 0;
      _tmp_284 <= 0;
      _tmp_285 <= 0;
      _tmp_286 <= 0;
      _tmp_287 <= 0;
      _tmp_288 <= 0;
      _tmp_289 <= 0;
      _tmp_290 <= 0;
      _tmp_291 <= 0;
      _tmp_292 <= 0;
      _tmp_293 <= 0;
      _tmp_294 <= 0;
      _tmp_295 <= 0;
      _tmp_296 <= 0;
      _tmp_297 <= 0;
      _tmp_298 <= 0;
      _tmp_299 <= 0;
      _tmp_300 <= 0;
      _tmp_301 <= 0;
      _tmp_302 <= 0;
      _tmp_303 <= 0;
      _tmp_304 <= 0;
      _tmp_305 <= 0;
      _tmp_306 <= 0;
      _tmp_307 <= 0;
      _tmp_308 <= 0;
      _tmp_309 <= 0;
      _tmp_310 <= 0;
      _tmp_311 <= 0;
      _tmp_312 <= 0;
      _tmp_313 <= 0;
      _tmp_314 <= 0;
      _tmp_315 <= 0;
      _tmp_316 <= 0;
      _tmp_317 <= 0;
      _tmp_318 <= 0;
      _tmp_319 <= 0;
      _tmp_320 <= 0;
      _tmp_321 <= 0;
      _tmp_322 <= 0;
      _tmp_323 <= 0;
      _tmp_324 <= 0;
      _tmp_325 <= 0;
      _tmp_326 <= 0;
      _tmp_327 <= 0;
      _tmp_328 <= 0;
      _tmp_329 <= 0;
      _tmp_330 <= 0;
      _tmp_331 <= 0;
      _tmp_332 <= 0;
      _tmp_333 <= 0;
      _tmp_334 <= 0;
      _tmp_335 <= 0;
      _tmp_336 <= 0;
      _tmp_337 <= 0;
      _tmp_338 <= 0;
      _tmp_339 <= 0;
      _tmp_340 <= 0;
      _tmp_341 <= 0;
      _tmp_342 <= 0;
      _tmp_343 <= 0;
      _tmp_344 <= 0;
      _tmp_345 <= 0;
      _stream_conv2d_2_sink_50_sink_mode <= 5'b0;
      _stream_conv2d_2_sink_50_sink_offset <= 0;
      _stream_conv2d_2_sink_50_sink_size <= 0;
      _stream_conv2d_2_sink_50_sink_stride <= 0;
      _stream_conv2d_2_sink_50_sink_sel <= 0;
      _stream_conv2d_2_sink_50_sink_offset_buf <= 0;
      _stream_conv2d_2_sink_50_sink_size_buf <= 0;
      _stream_conv2d_2_sink_50_sink_stride_buf <= 0;
      _stream_conv2d_2_sink_50_sink_waddr <= 0;
      _stream_conv2d_2_sink_50_sink_count <= 0;
      _stream_conv2d_2_sink_50_sink_wdata <= 0;
      _tmp_735 <= 0;
      _tmp_736 <= 0;
      _tmp_737 <= 0;
      _tmp_738 <= 0;
      _tmp_739 <= 0;
      _tmp_740 <= 0;
      __variable_wdata_264 <= 0;
      _tmp_741 <= 0;
      _tmp_742 <= 0;
      _tmp_743 <= 0;
      _tmp_744 <= 0;
      _tmp_747 <= 0;
      _tmp_750 <= 0;
      _tmp_751 <= 0;
      _tmp_752 <= 0;
      _tmp_753 <= 0;
      _tmp_754 <= 0;
      _tmp_755 <= 0;
      _tmp_756 <= 0;
      _tmp_757 <= 0;
      _tmp_758 <= 0;
      _tmp_759 <= 0;
      _tmp_760 <= 0;
      _tmp_761 <= 0;
      _tmp_762 <= 0;
      _tmp_763 <= 0;
      _tmp_764 <= 0;
      _tmp_765 <= 0;
      _tmp_766 <= 0;
      _tmp_767 <= 0;
      _tmp_768 <= 0;
      _tmp_769 <= 0;
      _tmp_770 <= 0;
      _tmp_771 <= 0;
      _tmp_772 <= 0;
      _tmp_773 <= 0;
      _tmp_774 <= 0;
      _tmp_775 <= 0;
      _tmp_776 <= 0;
      _tmp_777 <= 0;
      _tmp_778 <= 0;
      _tmp_779 <= 0;
      _tmp_780 <= 0;
      _tmp_781 <= 0;
      _tmp_782 <= 0;
      _tmp_783 <= 0;
      _tmp_784 <= 0;
      _tmp_785 <= 0;
      _tmp_786 <= 0;
      _tmp_787 <= 0;
      _tmp_788 <= 0;
      _tmp_789 <= 0;
      _tmp_790 <= 0;
      _tmp_791 <= 0;
      _tmp_792 <= 0;
      _tmp_793 <= 0;
      _tmp_794 <= 0;
      _tmp_795 <= 0;
      _tmp_796 <= 0;
      _tmp_797 <= 0;
      _tmp_798 <= 0;
      _tmp_799 <= 0;
      _tmp_800 <= 0;
      _tmp_801 <= 0;
      _tmp_802 <= 0;
      _tmp_803 <= 0;
      _tmp_804 <= 0;
      _tmp_805 <= 0;
      _tmp_806 <= 0;
      _tmp_807 <= 0;
      _tmp_808 <= 0;
      _tmp_809 <= 0;
      _tmp_810 <= 0;
      _tmp_811 <= 0;
      _tmp_812 <= 0;
      _tmp_813 <= 0;
      _tmp_814 <= 0;
      _tmp_815 <= 0;
      _tmp_816 <= 0;
      _tmp_817 <= 0;
      _tmp_818 <= 0;
      _tmp_819 <= 0;
      _tmp_820 <= 0;
      _tmp_821 <= 0;
      _tmp_822 <= 0;
      _tmp_823 <= 0;
      _tmp_824 <= 0;
      _tmp_825 <= 0;
      _tmp_826 <= 0;
      _tmp_827 <= 0;
      _tmp_828 <= 0;
      _tmp_829 <= 0;
      _tmp_830 <= 0;
      _tmp_831 <= 0;
      _tmp_832 <= 0;
      _tmp_833 <= 0;
      _tmp_834 <= 0;
      _tmp_835 <= 0;
      _tmp_836 <= 0;
      _tmp_837 <= 0;
      _tmp_838 <= 0;
      _tmp_839 <= 0;
      _tmp_840 <= 0;
      _tmp_841 <= 0;
      _tmp_842 <= 0;
      _tmp_843 <= 0;
      _tmp_844 <= 0;
      _stream_conv2d_2_busy_reg <= 0;
    end else begin
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_7_source_ram_renable <= 0;
        _stream_conv2d_2_source_7_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_7_idle <= _stream_conv2d_2_source_7_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_9_source_ram_renable <= 0;
        _stream_conv2d_2_source_9_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_9_idle <= _stream_conv2d_2_source_9_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_11_source_ram_renable <= 0;
        _stream_conv2d_2_source_11_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_11_idle <= _stream_conv2d_2_source_11_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_13_source_ram_renable <= 0;
        _stream_conv2d_2_source_13_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_13_idle <= _stream_conv2d_2_source_13_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_15_source_ram_renable <= 0;
        _stream_conv2d_2_source_15_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_15_idle <= _stream_conv2d_2_source_15_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_20_source_ram_renable <= 0;
        _stream_conv2d_2_source_20_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_20_idle <= _stream_conv2d_2_source_20_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_21_source_ram_renable <= 0;
        _stream_conv2d_2_source_21_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_21_idle <= _stream_conv2d_2_source_21_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_22_source_ram_renable <= 0;
        _stream_conv2d_2_source_22_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_22_idle <= _stream_conv2d_2_source_22_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_23_source_ram_renable <= 0;
        _stream_conv2d_2_source_23_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_23_idle <= _stream_conv2d_2_source_23_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_24_source_ram_renable <= 0;
        _stream_conv2d_2_source_24_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_24_idle <= _stream_conv2d_2_source_24_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_25_source_ram_renable <= 0;
        _stream_conv2d_2_source_25_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_25_idle <= _stream_conv2d_2_source_25_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_26_source_ram_renable <= 0;
        _stream_conv2d_2_source_26_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_26_idle <= _stream_conv2d_2_source_26_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_27_source_ram_renable <= 0;
        _stream_conv2d_2_source_27_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_27_idle <= _stream_conv2d_2_source_27_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_28_source_ram_renable <= 0;
        _stream_conv2d_2_source_28_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_28_idle <= _stream_conv2d_2_source_28_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_29_source_ram_renable <= 0;
        _stream_conv2d_2_source_29_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_29_idle <= _stream_conv2d_2_source_29_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_30_source_ram_renable <= 0;
        _stream_conv2d_2_source_30_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_30_idle <= _stream_conv2d_2_source_30_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_31_source_ram_renable <= 0;
        _stream_conv2d_2_source_31_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_31_idle <= _stream_conv2d_2_source_31_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_32_source_ram_renable <= 0;
        _stream_conv2d_2_source_32_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_32_idle <= _stream_conv2d_2_source_32_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_33_source_ram_renable <= 0;
        _stream_conv2d_2_source_33_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_33_idle <= _stream_conv2d_2_source_33_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_34_source_ram_renable <= 0;
        _stream_conv2d_2_source_34_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_34_idle <= _stream_conv2d_2_source_34_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_35_source_ram_renable <= 0;
        _stream_conv2d_2_source_35_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_35_idle <= _stream_conv2d_2_source_35_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_36_source_ram_renable <= 0;
        _stream_conv2d_2_source_36_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_36_idle <= _stream_conv2d_2_source_36_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_37_source_ram_renable <= 0;
        _stream_conv2d_2_source_37_source_fifo_deq <= 0;
      end 
      _stream_conv2d_2_source_37_idle <= _stream_conv2d_2_source_37_idle;
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_sink_50_sink_wenable <= 0;
        _stream_conv2d_2_sink_50_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_sink_51_sink_wenable <= 0;
        _stream_conv2d_2_sink_51_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_1 <= _stream_conv2d_2_stream_ivalid;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_2 <= __stream_conv2d_2_stream_ivalid_1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_3 <= __stream_conv2d_2_stream_ivalid_2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_4 <= __stream_conv2d_2_stream_ivalid_3;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_5 <= __stream_conv2d_2_stream_ivalid_4;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_6 <= __stream_conv2d_2_stream_ivalid_5;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_7 <= __stream_conv2d_2_stream_ivalid_6;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_8 <= __stream_conv2d_2_stream_ivalid_7;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_9 <= __stream_conv2d_2_stream_ivalid_8;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_10 <= __stream_conv2d_2_stream_ivalid_9;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_11 <= __stream_conv2d_2_stream_ivalid_10;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_12 <= __stream_conv2d_2_stream_ivalid_11;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_13 <= __stream_conv2d_2_stream_ivalid_12;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_14 <= __stream_conv2d_2_stream_ivalid_13;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_15 <= __stream_conv2d_2_stream_ivalid_14;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_16 <= __stream_conv2d_2_stream_ivalid_15;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_17 <= __stream_conv2d_2_stream_ivalid_16;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_18 <= __stream_conv2d_2_stream_ivalid_17;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_19 <= __stream_conv2d_2_stream_ivalid_18;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_20 <= __stream_conv2d_2_stream_ivalid_19;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_21 <= __stream_conv2d_2_stream_ivalid_20;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_22 <= __stream_conv2d_2_stream_ivalid_21;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_23 <= __stream_conv2d_2_stream_ivalid_22;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_24 <= __stream_conv2d_2_stream_ivalid_23;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_25 <= __stream_conv2d_2_stream_ivalid_24;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_26 <= __stream_conv2d_2_stream_ivalid_25;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_27 <= __stream_conv2d_2_stream_ivalid_26;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_28 <= __stream_conv2d_2_stream_ivalid_27;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __stream_conv2d_2_stream_ivalid_29 <= __stream_conv2d_2_stream_ivalid_28;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_322 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_326 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_329 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_332 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_336 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_339 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_342 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_346 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_349 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_352 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_356 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_359 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_362 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_366 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_369 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_372 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_376 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_379 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_382 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_386 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_389 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_392 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_396 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_399 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_402 <= stream_conv2d_2_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_406 <= stream_conv2d_2_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_409 <= stream_conv2d_2_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_412 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_416 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_419 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_422 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_426 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_429 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_432 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_436 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_439 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_442 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_446 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_449 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_452 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_456 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_459 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_462 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_466 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_469 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_472 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_476 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_479 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_482 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_486 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_489 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_492 <= stream_conv2d_2_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_496 <= stream_conv2d_2_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _eq_data_499 <= stream_conv2d_2_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_654 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_673 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_692 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_711 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_730 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_749 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_768 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_787 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_806 <= _cond_data_294 + stream_conv2d_2_parameter_16_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_822 <= _cond_data_301 + stream_conv2d_2_parameter_17_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_841 <= _cond_data_308 + stream_conv2d_2_parameter_18_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_866__variable_315 <= stream_conv2d_2_source_22_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_867__variable_314 <= stream_conv2d_2_source_21_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_868__variable_313 <= stream_conv2d_2_source_20_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_869__variable_318 <= stream_conv2d_2_source_25_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_870__variable_317 <= stream_conv2d_2_source_24_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_871__variable_316 <= stream_conv2d_2_source_23_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_872__variable_321 <= stream_conv2d_2_source_28_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_873__variable_320 <= stream_conv2d_2_source_27_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_874__variable_319 <= stream_conv2d_2_source_26_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_875_pointer_601 <= _pointer_data_601;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_876_reinterpretcast_592 <= _reinterpretcast_data_592;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_877_pointer_603 <= _pointer_data_603;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_878_reinterpretcast_593 <= _reinterpretcast_data_593;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_879_pointer_605 <= _pointer_data_605;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_880_reinterpretcast_594 <= _reinterpretcast_data_594;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_881_pointer_607 <= _pointer_data_607;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_882_reinterpretcast_595 <= _reinterpretcast_data_595;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_883_pointer_609 <= _pointer_data_609;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_884_reinterpretcast_596 <= _reinterpretcast_data_596;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_885_pointer_611 <= _pointer_data_611;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_886_reinterpretcast_597 <= _reinterpretcast_data_597;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_887_pointer_613 <= _pointer_data_613;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_888_reinterpretcast_598 <= _reinterpretcast_data_598;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_889_pointer_615 <= _pointer_data_615;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_890_reinterpretcast_599 <= _reinterpretcast_data_599;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_891_pointer_617 <= _pointer_data_617;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_892_reinterpretcast_600 <= _reinterpretcast_data_600;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_893__variable_264 <= stream_conv2d_2__reduce_reset_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_918__variable_259 <= stream_conv2d_2_parameter_0_data;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_931_cond_280 <= _cond_data_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_950_cond_287 <= _cond_data_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_894__delay_893__variable_264 <= __delay_data_893__variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_906_plus_822 <= _plus_data_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_919__delay_918__variable_259 <= __delay_data_918__variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_932__delay_931_cond_280 <= __delay_data_931_cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_951__delay_950_cond_287 <= __delay_data_950_cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_970_plus_841 <= _plus_data_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_895__delay_894__delay_893__variable_264 <= __delay_data_894__delay_893__variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_907__delay_906_plus_822 <= __delay_data_906_plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_920__delay_919__delay_918__variable_259 <= __delay_data_919__delay_918__variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_933__delay_932__delay_931_cond_280 <= __delay_data_932__delay_931_cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_952__delay_951__delay_950_cond_287 <= __delay_data_951__delay_950_cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_971__delay_970_plus_841 <= __delay_data_970_plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_896__delay_895__delay_894____variable_264 <= __delay_data_895__delay_894__delay_893__variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_908__delay_907__delay_906_plus_822 <= __delay_data_907__delay_906_plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_921__delay_920__delay_919____variable_259 <= __delay_data_920__delay_919__delay_918__variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_934__delay_933__delay_932__delay_931_cond_280 <= __delay_data_933__delay_932__delay_931_cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_953__delay_952__delay_951__delay_950_cond_287 <= __delay_data_952__delay_951__delay_950_cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_972__delay_971__delay_970_plus_841 <= __delay_data_971__delay_970_plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_897__delay_896__delay_895____variable_264 <= __delay_data_896__delay_895__delay_894____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_909__delay_908__delay_907__delay_906_plus_822 <= __delay_data_908__delay_907__delay_906_plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_922__delay_921__delay_920____variable_259 <= __delay_data_921__delay_920__delay_919____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_935__delay_934__delay_933__delay_932___cond_280 <= __delay_data_934__delay_933__delay_932__delay_931_cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_954__delay_953__delay_952__delay_951___cond_287 <= __delay_data_953__delay_952__delay_951__delay_950_cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_973__delay_972__delay_971__delay_970_plus_841 <= __delay_data_972__delay_971__delay_970_plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_898__delay_897__delay_896____variable_264 <= __delay_data_897__delay_896__delay_895____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_910__delay_909__delay_908__delay_907___plus_822 <= __delay_data_909__delay_908__delay_907__delay_906_plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_923__delay_922__delay_921____variable_259 <= __delay_data_922__delay_921__delay_920____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_936__delay_935__delay_934__delay_933___cond_280 <= __delay_data_935__delay_934__delay_933__delay_932___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_955__delay_954__delay_953__delay_952___cond_287 <= __delay_data_954__delay_953__delay_952__delay_951___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_974__delay_973__delay_972__delay_971___plus_841 <= __delay_data_973__delay_972__delay_971__delay_970_plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_899__delay_898__delay_897____variable_264 <= __delay_data_898__delay_897__delay_896____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_911__delay_910__delay_909__delay_908___plus_822 <= __delay_data_910__delay_909__delay_908__delay_907___plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_924__delay_923__delay_922____variable_259 <= __delay_data_923__delay_922__delay_921____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_937__delay_936__delay_935__delay_934___cond_280 <= __delay_data_936__delay_935__delay_934__delay_933___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_956__delay_955__delay_954__delay_953___cond_287 <= __delay_data_955__delay_954__delay_953__delay_952___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_975__delay_974__delay_973__delay_972___plus_841 <= __delay_data_974__delay_973__delay_972__delay_971___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_900__delay_899__delay_898____variable_264 <= __delay_data_899__delay_898__delay_897____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_912__delay_911__delay_910__delay_909___plus_822 <= __delay_data_911__delay_910__delay_909__delay_908___plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_925__delay_924__delay_923____variable_259 <= __delay_data_924__delay_923__delay_922____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_938__delay_937__delay_936__delay_935___cond_280 <= __delay_data_937__delay_936__delay_935__delay_934___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_957__delay_956__delay_955__delay_954___cond_287 <= __delay_data_956__delay_955__delay_954__delay_953___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_976__delay_975__delay_974__delay_973___plus_841 <= __delay_data_975__delay_974__delay_973__delay_972___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_901__delay_900__delay_899____variable_264 <= __delay_data_900__delay_899__delay_898____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_913__delay_912__delay_911__delay_910___plus_822 <= __delay_data_912__delay_911__delay_910__delay_909___plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_926__delay_925__delay_924____variable_259 <= __delay_data_925__delay_924__delay_923____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_939__delay_938__delay_937__delay_936___cond_280 <= __delay_data_938__delay_937__delay_936__delay_935___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_958__delay_957__delay_956__delay_955___cond_287 <= __delay_data_957__delay_956__delay_955__delay_954___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_977__delay_976__delay_975__delay_974___plus_841 <= __delay_data_976__delay_975__delay_974__delay_973___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_902__delay_901__delay_900____variable_264 <= __delay_data_901__delay_900__delay_899____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_914__delay_913__delay_912__delay_911___plus_822 <= __delay_data_913__delay_912__delay_911__delay_910___plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_927__delay_926__delay_925____variable_259 <= __delay_data_926__delay_925__delay_924____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_940__delay_939__delay_938__delay_937___cond_280 <= __delay_data_939__delay_938__delay_937__delay_936___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_959__delay_958__delay_957__delay_956___cond_287 <= __delay_data_958__delay_957__delay_956__delay_955___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_978__delay_977__delay_976__delay_975___plus_841 <= __delay_data_977__delay_976__delay_975__delay_974___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_903__delay_902__delay_901____variable_264 <= __delay_data_902__delay_901__delay_900____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_915__delay_914__delay_913__delay_912___plus_822 <= __delay_data_914__delay_913__delay_912__delay_911___plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_928__delay_927__delay_926____variable_259 <= __delay_data_927__delay_926__delay_925____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_941__delay_940__delay_939__delay_938___cond_280 <= __delay_data_940__delay_939__delay_938__delay_937___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_960__delay_959__delay_958__delay_957___cond_287 <= __delay_data_959__delay_958__delay_957__delay_956___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_979__delay_978__delay_977__delay_976___plus_841 <= __delay_data_978__delay_977__delay_976__delay_975___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_904__delay_903__delay_902____variable_264 <= __delay_data_903__delay_902__delay_901____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_916__delay_915__delay_914__delay_913___plus_822 <= __delay_data_915__delay_914__delay_913__delay_912___plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_929__delay_928__delay_927____variable_259 <= __delay_data_928__delay_927__delay_926____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_942__delay_941__delay_940__delay_939___cond_280 <= __delay_data_941__delay_940__delay_939__delay_938___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_961__delay_960__delay_959__delay_958___cond_287 <= __delay_data_960__delay_959__delay_958__delay_957___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_980__delay_979__delay_978__delay_977___plus_841 <= __delay_data_979__delay_978__delay_977__delay_976___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_905__delay_904__delay_903____variable_264 <= __delay_data_904__delay_903__delay_902____variable_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_917__delay_916__delay_915__delay_914___plus_822 <= __delay_data_916__delay_915__delay_914__delay_913___plus_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_930__delay_929__delay_928____variable_259 <= __delay_data_929__delay_928__delay_927____variable_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_943__delay_942__delay_941__delay_940___cond_280 <= __delay_data_942__delay_941__delay_940__delay_939___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_962__delay_961__delay_960__delay_959___cond_287 <= __delay_data_961__delay_960__delay_959__delay_958___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_981__delay_980__delay_979__delay_978___plus_841 <= __delay_data_980__delay_979__delay_978__delay_977___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_944__delay_943__delay_942__delay_941___cond_280 <= __delay_data_943__delay_942__delay_941__delay_940___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_963__delay_962__delay_961__delay_960___cond_287 <= __delay_data_962__delay_961__delay_960__delay_959___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_982__delay_981__delay_980__delay_979___plus_841 <= __delay_data_981__delay_980__delay_979__delay_978___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_945__delay_944__delay_943__delay_942___cond_280 <= __delay_data_944__delay_943__delay_942__delay_941___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_964__delay_963__delay_962__delay_961___cond_287 <= __delay_data_963__delay_962__delay_961__delay_960___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_983__delay_982__delay_981__delay_980___plus_841 <= __delay_data_982__delay_981__delay_980__delay_979___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_946__delay_945__delay_944__delay_943___cond_280 <= __delay_data_945__delay_944__delay_943__delay_942___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_965__delay_964__delay_963__delay_962___cond_287 <= __delay_data_964__delay_963__delay_962__delay_961___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_984__delay_983__delay_982__delay_981___plus_841 <= __delay_data_983__delay_982__delay_981__delay_980___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_947__delay_946__delay_945__delay_944___cond_280 <= __delay_data_946__delay_945__delay_944__delay_943___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_966__delay_965__delay_964__delay_963___cond_287 <= __delay_data_965__delay_964__delay_963__delay_962___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_985__delay_984__delay_983__delay_982___plus_841 <= __delay_data_984__delay_983__delay_982__delay_981___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_948__delay_947__delay_946__delay_945___cond_280 <= __delay_data_947__delay_946__delay_945__delay_944___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_967__delay_966__delay_965__delay_964___cond_287 <= __delay_data_966__delay_965__delay_964__delay_963___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_986__delay_985__delay_984__delay_983___plus_841 <= __delay_data_985__delay_984__delay_983__delay_982___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_949__delay_948__delay_947__delay_946___cond_280 <= __delay_data_948__delay_947__delay_946__delay_945___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_968__delay_967__delay_966__delay_965___cond_287 <= __delay_data_967__delay_966__delay_965__delay_964___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_987__delay_986__delay_985__delay_984___plus_841 <= __delay_data_986__delay_985__delay_984__delay_983___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _plus_data_825 <= __substreamoutput_data_823 + __delay_data_949__delay_948__delay_947__delay_946___cond_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_969__delay_968__delay_967__delay_966___cond_287 <= __delay_data_968__delay_967__delay_966__delay_965___cond_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_988__delay_987__delay_986__delay_985___plus_841 <= __delay_data_987__delay_986__delay_985__delay_984___plus_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_989__substreamoutput_824 <= __substreamoutput_data_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_990__delay_989__substreamoutput_824 <= __delay_data_989__substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_991__delay_990__delay_989__substreamoutput_824 <= __delay_data_990__delay_989__substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_992__delay_991__delay_990____substreamoutput_824 <= __delay_data_991__delay_990__delay_989__substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_993__delay_992__delay_991____substreamoutput_824 <= __delay_data_992__delay_991__delay_990____substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_994__delay_993__delay_992____substreamoutput_824 <= __delay_data_993__delay_992__delay_991____substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_995__delay_994__delay_993____substreamoutput_824 <= __delay_data_994__delay_993__delay_992____substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_996__delay_995__delay_994____substreamoutput_824 <= __delay_data_995__delay_994__delay_993____substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_997__delay_996__delay_995____substreamoutput_824 <= __delay_data_996__delay_995__delay_994____substreamoutput_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        __delay_data_998__delay_997__delay_996____substreamoutput_824 <= __delay_data_997__delay_996__delay_995____substreamoutput_824;
      end 
      if(_set_flag_177) begin
        _stream_conv2d_2_parameter_0_next_parameter_data <= cparam_conv2d_2_stream_reduce_size;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_259 <= _stream_conv2d_2_parameter_0_next_parameter_data;
      end 
      if(_set_flag_178) begin
        _stream_conv2d_2_parameter_1_next_parameter_data <= conv2d_2_col_select;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_260 <= _stream_conv2d_2_parameter_1_next_parameter_data;
      end 
      if(_set_flag_179) begin
        _stream_conv2d_2_parameter_2_next_parameter_data <= conv2d_2_row_select_buf;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_261 <= _stream_conv2d_2_parameter_2_next_parameter_data;
      end 
      if(_set_flag_180) begin
        _stream_conv2d_2_parameter_3_next_parameter_data <= conv2d_2_stream_pad_masks;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_262 <= _stream_conv2d_2_parameter_3_next_parameter_data;
      end 
      if(_set_flag_181) begin
        _stream_conv2d_2_parameter_4_next_parameter_data <= cparam_conv2d_2_stream_omit_mask;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_263 <= _stream_conv2d_2_parameter_4_next_parameter_data;
      end 
      if(_set_flag_182) begin
        _stream_conv2d_2_parameter_6_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_274 <= _stream_conv2d_2_parameter_6_next_parameter_data;
      end 
      if(_set_flag_183) begin
        _stream_conv2d_2_source_7_source_mode <= 5'b0;
        _stream_conv2d_2_source_7_source_empty_data <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_7_source_mode & 5'b0))) begin
        _stream_conv2d_2_source_7_idle <= 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_7_source_mode & 5'b0)) && _stream_conv2d_2_is_root) begin
        __variable_wdata_275 <= _stream_conv2d_2_source_7_source_empty_data;
      end 
      if(_set_flag_184) begin
        _stream_conv2d_2_parameter_8_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_281 <= _stream_conv2d_2_parameter_8_next_parameter_data;
      end 
      if(_set_flag_185) begin
        _stream_conv2d_2_source_9_source_mode <= 5'b0;
        _stream_conv2d_2_source_9_source_empty_data <= 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_9_source_mode & 5'b0))) begin
        _stream_conv2d_2_source_9_idle <= 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_9_source_mode & 5'b0)) && _stream_conv2d_2_is_root) begin
        __variable_wdata_282 <= _stream_conv2d_2_source_9_source_empty_data;
      end 
      if(_set_flag_186) begin
        _stream_conv2d_2_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_288 <= _stream_conv2d_2_parameter_10_next_parameter_data;
      end 
      if(_set_flag_187) begin
        _stream_conv2d_2_source_11_source_mode <= 5'b0;
        _stream_conv2d_2_source_11_source_empty_data <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_11_source_mode & 5'b0))) begin
        _stream_conv2d_2_source_11_idle <= 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_11_source_mode & 5'b0)) && _stream_conv2d_2_is_root) begin
        __variable_wdata_289 <= _stream_conv2d_2_source_11_source_empty_data;
      end 
      if(_set_flag_188) begin
        _stream_conv2d_2_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_295 <= _stream_conv2d_2_parameter_12_next_parameter_data;
      end 
      if(_set_flag_189) begin
        _stream_conv2d_2_source_13_source_mode <= 5'b0;
        _stream_conv2d_2_source_13_source_empty_data <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_13_source_mode & 5'b0))) begin
        _stream_conv2d_2_source_13_idle <= 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_13_source_mode & 5'b0)) && _stream_conv2d_2_is_root) begin
        __variable_wdata_296 <= _stream_conv2d_2_source_13_source_empty_data;
      end 
      if(_set_flag_190) begin
        _stream_conv2d_2_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_302 <= _stream_conv2d_2_parameter_14_next_parameter_data;
      end 
      if(_set_flag_191) begin
        _stream_conv2d_2_source_15_source_mode <= 5'b0;
        _stream_conv2d_2_source_15_source_empty_data <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_15_source_mode & 5'b0))) begin
        _stream_conv2d_2_source_15_idle <= 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready && !(|(_stream_conv2d_2_source_15_source_mode & 5'b0)) && _stream_conv2d_2_is_root) begin
        __variable_wdata_303 <= _stream_conv2d_2_source_15_source_empty_data;
      end 
      if(_set_flag_192) begin
        _stream_conv2d_2_parameter_16_next_parameter_data <= cparam_conv2d_2_cshamt_mul_value;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_309 <= _stream_conv2d_2_parameter_16_next_parameter_data;
      end 
      if(_set_flag_193) begin
        _stream_conv2d_2_parameter_17_next_parameter_data <= cparam_conv2d_2_cshamt_sum_value;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_310 <= _stream_conv2d_2_parameter_17_next_parameter_data;
      end 
      if(_set_flag_194) begin
        _stream_conv2d_2_parameter_18_next_parameter_data <= cparam_conv2d_2_cshamt_out_value;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_311 <= _stream_conv2d_2_parameter_18_next_parameter_data;
      end 
      if(_set_flag_195) begin
        _stream_conv2d_2_parameter_19_next_parameter_data <= cparam_conv2d_2_act_func_index;
      end 
      if(_stream_conv2d_2_source_start) begin
        __variable_wdata_312 <= _stream_conv2d_2_parameter_19_next_parameter_data;
      end 
      if(_set_flag_196) begin
        _stream_conv2d_2_source_20_source_mode <= 5'b10;
        _stream_conv2d_2_source_20_source_offset <= conv2d_2_stream_act_local_0 + conv2d_2_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_196) begin
        _source_stream_conv2d_2_source_20_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_196) begin
        _source_stream_conv2d_2_source_20_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_196) begin
        _source_stream_conv2d_2_source_20_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_196) begin
        _source_stream_conv2d_2_source_20_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_196) begin
        _stream_conv2d_2_source_20_source_sel <= 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_20_source_offset_buf <= _stream_conv2d_2_source_20_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_count_0 <= _source_stream_conv2d_2_source_20_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_count_1 <= _source_stream_conv2d_2_source_20_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_count_2 <= _source_stream_conv2d_2_source_20_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_count_3 <= _source_stream_conv2d_2_source_20_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_size_buf_0 <= _source_stream_conv2d_2_source_20_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_size_buf_1 <= _source_stream_conv2d_2_source_20_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_size_buf_2 <= _source_stream_conv2d_2_source_20_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_size_buf_3 <= _source_stream_conv2d_2_source_20_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_stride_buf_0 <= _source_stream_conv2d_2_source_20_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_stride_buf_1 <= _source_stream_conv2d_2_source_20_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_stride_buf_2 <= _source_stream_conv2d_2_source_20_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_stride_buf_3 <= _source_stream_conv2d_2_source_20_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_313 <= _stream_conv2d_2_source_20_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_20_idle <= 0;
        _stream_conv2d_2_source_20_source_ram_raddr <= _stream_conv2d_2_source_20_source_pat_all_offset;
        _stream_conv2d_2_source_20_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_0 <= _source_stream_conv2d_2_source_20_pat_cur_offset_0 + _source_stream_conv2d_2_source_20_pat_stride_buf_0;
        _source_stream_conv2d_2_source_20_pat_count_0 <= _source_stream_conv2d_2_source_20_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && (_source_stream_conv2d_2_source_20_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_20_pat_count_0 <= _source_stream_conv2d_2_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && (_source_stream_conv2d_2_source_20_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_1 <= _source_stream_conv2d_2_source_20_pat_cur_offset_1 + _source_stream_conv2d_2_source_20_pat_stride_buf_1;
        _source_stream_conv2d_2_source_20_pat_count_1 <= _source_stream_conv2d_2_source_20_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && (_source_stream_conv2d_2_source_20_pat_count_0 == 0) && (_source_stream_conv2d_2_source_20_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_20_pat_count_1 <= _source_stream_conv2d_2_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_2_source_20_pat_count_0 == 0) && (_source_stream_conv2d_2_source_20_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_2 <= _source_stream_conv2d_2_source_20_pat_cur_offset_2 + _source_stream_conv2d_2_source_20_pat_stride_buf_2;
        _source_stream_conv2d_2_source_20_pat_count_2 <= _source_stream_conv2d_2_source_20_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_2_source_20_pat_count_0 == 0) && (_source_stream_conv2d_2_source_20_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_20_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_20_pat_count_2 <= _source_stream_conv2d_2_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_2_source_20_pat_count_0 == 0) && (_source_stream_conv2d_2_source_20_pat_count_1 == 0) && (_source_stream_conv2d_2_source_20_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_3 <= _source_stream_conv2d_2_source_20_pat_cur_offset_3 + _source_stream_conv2d_2_source_20_pat_stride_buf_3;
        _source_stream_conv2d_2_source_20_pat_count_3 <= _source_stream_conv2d_2_source_20_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_2_source_20_pat_count_0 == 0) && (_source_stream_conv2d_2_source_20_pat_count_1 == 0) && (_source_stream_conv2d_2_source_20_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_20_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_20_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_20_pat_count_3 <= _source_stream_conv2d_2_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_20_source_ram_renable <= 0;
        _stream_conv2d_2_source_20_idle <= 1;
      end 
      if((_stream_conv2d_2_source_20_source_pat_fsm_0 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_20_source_ram_renable <= 0;
        _stream_conv2d_2_source_20_idle <= 1;
      end 
      if(_set_flag_199) begin
        _stream_conv2d_2_source_21_source_mode <= 5'b10;
        _stream_conv2d_2_source_21_source_offset <= conv2d_2_stream_act_local_1 + conv2d_2_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_199) begin
        _source_stream_conv2d_2_source_21_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_199) begin
        _source_stream_conv2d_2_source_21_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_21_pat_stride_1 <= 0;
      end 
      if(_set_flag_199) begin
        _source_stream_conv2d_2_source_21_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_199) begin
        _source_stream_conv2d_2_source_21_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_199) begin
        _stream_conv2d_2_source_21_source_sel <= 2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_21_source_offset_buf <= _stream_conv2d_2_source_21_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_count_0 <= _source_stream_conv2d_2_source_21_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_count_1 <= _source_stream_conv2d_2_source_21_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_count_2 <= _source_stream_conv2d_2_source_21_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_count_3 <= _source_stream_conv2d_2_source_21_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_size_buf_0 <= _source_stream_conv2d_2_source_21_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_size_buf_1 <= _source_stream_conv2d_2_source_21_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_size_buf_2 <= _source_stream_conv2d_2_source_21_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_size_buf_3 <= _source_stream_conv2d_2_source_21_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_stride_buf_0 <= _source_stream_conv2d_2_source_21_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_stride_buf_1 <= _source_stream_conv2d_2_source_21_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_stride_buf_2 <= _source_stream_conv2d_2_source_21_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_stride_buf_3 <= _source_stream_conv2d_2_source_21_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_314 <= _stream_conv2d_2_source_21_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_21_idle <= 0;
        _stream_conv2d_2_source_21_source_ram_raddr <= _stream_conv2d_2_source_21_source_pat_all_offset;
        _stream_conv2d_2_source_21_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_0 <= _source_stream_conv2d_2_source_21_pat_cur_offset_0 + _source_stream_conv2d_2_source_21_pat_stride_buf_0;
        _source_stream_conv2d_2_source_21_pat_count_0 <= _source_stream_conv2d_2_source_21_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && (_source_stream_conv2d_2_source_21_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_21_pat_count_0 <= _source_stream_conv2d_2_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && (_source_stream_conv2d_2_source_21_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_1 <= _source_stream_conv2d_2_source_21_pat_cur_offset_1 + _source_stream_conv2d_2_source_21_pat_stride_buf_1;
        _source_stream_conv2d_2_source_21_pat_count_1 <= _source_stream_conv2d_2_source_21_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && (_source_stream_conv2d_2_source_21_pat_count_0 == 0) && (_source_stream_conv2d_2_source_21_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_21_pat_count_1 <= _source_stream_conv2d_2_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_2_source_21_pat_count_0 == 0) && (_source_stream_conv2d_2_source_21_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_2 <= _source_stream_conv2d_2_source_21_pat_cur_offset_2 + _source_stream_conv2d_2_source_21_pat_stride_buf_2;
        _source_stream_conv2d_2_source_21_pat_count_2 <= _source_stream_conv2d_2_source_21_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_2_source_21_pat_count_0 == 0) && (_source_stream_conv2d_2_source_21_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_21_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_21_pat_count_2 <= _source_stream_conv2d_2_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_2_source_21_pat_count_0 == 0) && (_source_stream_conv2d_2_source_21_pat_count_1 == 0) && (_source_stream_conv2d_2_source_21_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_3 <= _source_stream_conv2d_2_source_21_pat_cur_offset_3 + _source_stream_conv2d_2_source_21_pat_stride_buf_3;
        _source_stream_conv2d_2_source_21_pat_count_3 <= _source_stream_conv2d_2_source_21_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_2_source_21_pat_count_0 == 0) && (_source_stream_conv2d_2_source_21_pat_count_1 == 0) && (_source_stream_conv2d_2_source_21_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_21_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_21_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_21_pat_count_3 <= _source_stream_conv2d_2_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_21_source_ram_renable <= 0;
        _stream_conv2d_2_source_21_idle <= 1;
      end 
      if((_stream_conv2d_2_source_21_source_pat_fsm_1 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_21_source_ram_renable <= 0;
        _stream_conv2d_2_source_21_idle <= 1;
      end 
      if(_set_flag_202) begin
        _stream_conv2d_2_source_22_source_mode <= 5'b10;
        _stream_conv2d_2_source_22_source_offset <= conv2d_2_stream_act_local_2 + conv2d_2_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_202) begin
        _source_stream_conv2d_2_source_22_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_202) begin
        _source_stream_conv2d_2_source_22_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_22_pat_stride_1 <= 0;
      end 
      if(_set_flag_202) begin
        _source_stream_conv2d_2_source_22_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_202) begin
        _source_stream_conv2d_2_source_22_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_202) begin
        _stream_conv2d_2_source_22_source_sel <= 3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_22_source_offset_buf <= _stream_conv2d_2_source_22_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_count_0 <= _source_stream_conv2d_2_source_22_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_count_1 <= _source_stream_conv2d_2_source_22_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_count_2 <= _source_stream_conv2d_2_source_22_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_count_3 <= _source_stream_conv2d_2_source_22_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_size_buf_0 <= _source_stream_conv2d_2_source_22_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_size_buf_1 <= _source_stream_conv2d_2_source_22_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_size_buf_2 <= _source_stream_conv2d_2_source_22_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_size_buf_3 <= _source_stream_conv2d_2_source_22_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_stride_buf_0 <= _source_stream_conv2d_2_source_22_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_stride_buf_1 <= _source_stream_conv2d_2_source_22_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_stride_buf_2 <= _source_stream_conv2d_2_source_22_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_stride_buf_3 <= _source_stream_conv2d_2_source_22_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_315 <= _stream_conv2d_2_source_22_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_22_idle <= 0;
        _stream_conv2d_2_source_22_source_ram_raddr <= _stream_conv2d_2_source_22_source_pat_all_offset;
        _stream_conv2d_2_source_22_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_0 <= _source_stream_conv2d_2_source_22_pat_cur_offset_0 + _source_stream_conv2d_2_source_22_pat_stride_buf_0;
        _source_stream_conv2d_2_source_22_pat_count_0 <= _source_stream_conv2d_2_source_22_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && (_source_stream_conv2d_2_source_22_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_22_pat_count_0 <= _source_stream_conv2d_2_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && (_source_stream_conv2d_2_source_22_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_1 <= _source_stream_conv2d_2_source_22_pat_cur_offset_1 + _source_stream_conv2d_2_source_22_pat_stride_buf_1;
        _source_stream_conv2d_2_source_22_pat_count_1 <= _source_stream_conv2d_2_source_22_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && (_source_stream_conv2d_2_source_22_pat_count_0 == 0) && (_source_stream_conv2d_2_source_22_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_22_pat_count_1 <= _source_stream_conv2d_2_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_2_source_22_pat_count_0 == 0) && (_source_stream_conv2d_2_source_22_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_2 <= _source_stream_conv2d_2_source_22_pat_cur_offset_2 + _source_stream_conv2d_2_source_22_pat_stride_buf_2;
        _source_stream_conv2d_2_source_22_pat_count_2 <= _source_stream_conv2d_2_source_22_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_2_source_22_pat_count_0 == 0) && (_source_stream_conv2d_2_source_22_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_22_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_22_pat_count_2 <= _source_stream_conv2d_2_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_2_source_22_pat_count_0 == 0) && (_source_stream_conv2d_2_source_22_pat_count_1 == 0) && (_source_stream_conv2d_2_source_22_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_3 <= _source_stream_conv2d_2_source_22_pat_cur_offset_3 + _source_stream_conv2d_2_source_22_pat_stride_buf_3;
        _source_stream_conv2d_2_source_22_pat_count_3 <= _source_stream_conv2d_2_source_22_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_2_source_22_pat_count_0 == 0) && (_source_stream_conv2d_2_source_22_pat_count_1 == 0) && (_source_stream_conv2d_2_source_22_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_22_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_22_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_22_pat_count_3 <= _source_stream_conv2d_2_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_22_source_ram_renable <= 0;
        _stream_conv2d_2_source_22_idle <= 1;
      end 
      if((_stream_conv2d_2_source_22_source_pat_fsm_2 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_22_source_ram_renable <= 0;
        _stream_conv2d_2_source_22_idle <= 1;
      end 
      if(_set_flag_205) begin
        _stream_conv2d_2_source_23_source_mode <= 5'b10;
        _stream_conv2d_2_source_23_source_offset <= conv2d_2_stream_act_local_3 + conv2d_2_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_205) begin
        _source_stream_conv2d_2_source_23_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_23_pat_stride_0 <= 1;
      end 
      if(_set_flag_205) begin
        _source_stream_conv2d_2_source_23_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_23_pat_stride_1 <= 0;
      end 
      if(_set_flag_205) begin
        _source_stream_conv2d_2_source_23_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_23_pat_stride_2 <= 0;
      end 
      if(_set_flag_205) begin
        _source_stream_conv2d_2_source_23_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_23_pat_stride_3 <= 0;
      end 
      if(_set_flag_205) begin
        _stream_conv2d_2_source_23_source_sel <= 4;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_23_source_offset_buf <= _stream_conv2d_2_source_23_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_count_0 <= _source_stream_conv2d_2_source_23_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_count_1 <= _source_stream_conv2d_2_source_23_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_count_2 <= _source_stream_conv2d_2_source_23_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_count_3 <= _source_stream_conv2d_2_source_23_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_size_buf_0 <= _source_stream_conv2d_2_source_23_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_size_buf_1 <= _source_stream_conv2d_2_source_23_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_size_buf_2 <= _source_stream_conv2d_2_source_23_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_size_buf_3 <= _source_stream_conv2d_2_source_23_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_stride_buf_0 <= _source_stream_conv2d_2_source_23_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_stride_buf_1 <= _source_stream_conv2d_2_source_23_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_stride_buf_2 <= _source_stream_conv2d_2_source_23_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_stride_buf_3 <= _source_stream_conv2d_2_source_23_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_316 <= _stream_conv2d_2_source_23_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_23_idle <= 0;
        _stream_conv2d_2_source_23_source_ram_raddr <= _stream_conv2d_2_source_23_source_pat_all_offset;
        _stream_conv2d_2_source_23_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_0 <= _source_stream_conv2d_2_source_23_pat_cur_offset_0 + _source_stream_conv2d_2_source_23_pat_stride_buf_0;
        _source_stream_conv2d_2_source_23_pat_count_0 <= _source_stream_conv2d_2_source_23_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && (_source_stream_conv2d_2_source_23_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_23_pat_count_0 <= _source_stream_conv2d_2_source_23_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && (_source_stream_conv2d_2_source_23_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_1 <= _source_stream_conv2d_2_source_23_pat_cur_offset_1 + _source_stream_conv2d_2_source_23_pat_stride_buf_1;
        _source_stream_conv2d_2_source_23_pat_count_1 <= _source_stream_conv2d_2_source_23_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && (_source_stream_conv2d_2_source_23_pat_count_0 == 0) && (_source_stream_conv2d_2_source_23_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_23_pat_count_1 <= _source_stream_conv2d_2_source_23_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_2_source_23_pat_count_0 == 0) && (_source_stream_conv2d_2_source_23_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_2 <= _source_stream_conv2d_2_source_23_pat_cur_offset_2 + _source_stream_conv2d_2_source_23_pat_stride_buf_2;
        _source_stream_conv2d_2_source_23_pat_count_2 <= _source_stream_conv2d_2_source_23_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_2_source_23_pat_count_0 == 0) && (_source_stream_conv2d_2_source_23_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_23_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_23_pat_count_2 <= _source_stream_conv2d_2_source_23_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_2_source_23_pat_count_0 == 0) && (_source_stream_conv2d_2_source_23_pat_count_1 == 0) && (_source_stream_conv2d_2_source_23_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_3 <= _source_stream_conv2d_2_source_23_pat_cur_offset_3 + _source_stream_conv2d_2_source_23_pat_stride_buf_3;
        _source_stream_conv2d_2_source_23_pat_count_3 <= _source_stream_conv2d_2_source_23_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_2_source_23_pat_count_0 == 0) && (_source_stream_conv2d_2_source_23_pat_count_1 == 0) && (_source_stream_conv2d_2_source_23_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_23_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_23_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_23_pat_count_3 <= _source_stream_conv2d_2_source_23_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_23_source_ram_renable <= 0;
        _stream_conv2d_2_source_23_idle <= 1;
      end 
      if((_stream_conv2d_2_source_23_source_pat_fsm_3 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_23_source_ram_renable <= 0;
        _stream_conv2d_2_source_23_idle <= 1;
      end 
      if(_set_flag_208) begin
        _stream_conv2d_2_source_24_source_mode <= 5'b10;
        _stream_conv2d_2_source_24_source_offset <= conv2d_2_stream_act_local_4 + conv2d_2_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_208) begin
        _source_stream_conv2d_2_source_24_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_24_pat_stride_0 <= 1;
      end 
      if(_set_flag_208) begin
        _source_stream_conv2d_2_source_24_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_24_pat_stride_1 <= 0;
      end 
      if(_set_flag_208) begin
        _source_stream_conv2d_2_source_24_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_24_pat_stride_2 <= 0;
      end 
      if(_set_flag_208) begin
        _source_stream_conv2d_2_source_24_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_24_pat_stride_3 <= 0;
      end 
      if(_set_flag_208) begin
        _stream_conv2d_2_source_24_source_sel <= 5;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_24_source_offset_buf <= _stream_conv2d_2_source_24_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_count_0 <= _source_stream_conv2d_2_source_24_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_count_1 <= _source_stream_conv2d_2_source_24_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_count_2 <= _source_stream_conv2d_2_source_24_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_count_3 <= _source_stream_conv2d_2_source_24_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_size_buf_0 <= _source_stream_conv2d_2_source_24_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_size_buf_1 <= _source_stream_conv2d_2_source_24_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_size_buf_2 <= _source_stream_conv2d_2_source_24_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_size_buf_3 <= _source_stream_conv2d_2_source_24_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_stride_buf_0 <= _source_stream_conv2d_2_source_24_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_stride_buf_1 <= _source_stream_conv2d_2_source_24_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_stride_buf_2 <= _source_stream_conv2d_2_source_24_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_stride_buf_3 <= _source_stream_conv2d_2_source_24_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_317 <= _stream_conv2d_2_source_24_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_24_idle <= 0;
        _stream_conv2d_2_source_24_source_ram_raddr <= _stream_conv2d_2_source_24_source_pat_all_offset;
        _stream_conv2d_2_source_24_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_0 <= _source_stream_conv2d_2_source_24_pat_cur_offset_0 + _source_stream_conv2d_2_source_24_pat_stride_buf_0;
        _source_stream_conv2d_2_source_24_pat_count_0 <= _source_stream_conv2d_2_source_24_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && (_source_stream_conv2d_2_source_24_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_24_pat_count_0 <= _source_stream_conv2d_2_source_24_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && (_source_stream_conv2d_2_source_24_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_1 <= _source_stream_conv2d_2_source_24_pat_cur_offset_1 + _source_stream_conv2d_2_source_24_pat_stride_buf_1;
        _source_stream_conv2d_2_source_24_pat_count_1 <= _source_stream_conv2d_2_source_24_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && (_source_stream_conv2d_2_source_24_pat_count_0 == 0) && (_source_stream_conv2d_2_source_24_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_24_pat_count_1 <= _source_stream_conv2d_2_source_24_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_2_source_24_pat_count_0 == 0) && (_source_stream_conv2d_2_source_24_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_2 <= _source_stream_conv2d_2_source_24_pat_cur_offset_2 + _source_stream_conv2d_2_source_24_pat_stride_buf_2;
        _source_stream_conv2d_2_source_24_pat_count_2 <= _source_stream_conv2d_2_source_24_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_2_source_24_pat_count_0 == 0) && (_source_stream_conv2d_2_source_24_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_24_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_24_pat_count_2 <= _source_stream_conv2d_2_source_24_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_2_source_24_pat_count_0 == 0) && (_source_stream_conv2d_2_source_24_pat_count_1 == 0) && (_source_stream_conv2d_2_source_24_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_3 <= _source_stream_conv2d_2_source_24_pat_cur_offset_3 + _source_stream_conv2d_2_source_24_pat_stride_buf_3;
        _source_stream_conv2d_2_source_24_pat_count_3 <= _source_stream_conv2d_2_source_24_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_2_source_24_pat_count_0 == 0) && (_source_stream_conv2d_2_source_24_pat_count_1 == 0) && (_source_stream_conv2d_2_source_24_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_24_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_24_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_24_pat_count_3 <= _source_stream_conv2d_2_source_24_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_24_source_ram_renable <= 0;
        _stream_conv2d_2_source_24_idle <= 1;
      end 
      if((_stream_conv2d_2_source_24_source_pat_fsm_4 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_24_source_ram_renable <= 0;
        _stream_conv2d_2_source_24_idle <= 1;
      end 
      if(_set_flag_211) begin
        _stream_conv2d_2_source_25_source_mode <= 5'b10;
        _stream_conv2d_2_source_25_source_offset <= conv2d_2_stream_act_local_5 + conv2d_2_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_211) begin
        _source_stream_conv2d_2_source_25_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_25_pat_stride_0 <= 1;
      end 
      if(_set_flag_211) begin
        _source_stream_conv2d_2_source_25_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_25_pat_stride_1 <= 0;
      end 
      if(_set_flag_211) begin
        _source_stream_conv2d_2_source_25_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_25_pat_stride_2 <= 0;
      end 
      if(_set_flag_211) begin
        _source_stream_conv2d_2_source_25_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_25_pat_stride_3 <= 0;
      end 
      if(_set_flag_211) begin
        _stream_conv2d_2_source_25_source_sel <= 6;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_25_source_offset_buf <= _stream_conv2d_2_source_25_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_count_0 <= _source_stream_conv2d_2_source_25_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_count_1 <= _source_stream_conv2d_2_source_25_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_count_2 <= _source_stream_conv2d_2_source_25_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_count_3 <= _source_stream_conv2d_2_source_25_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_size_buf_0 <= _source_stream_conv2d_2_source_25_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_size_buf_1 <= _source_stream_conv2d_2_source_25_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_size_buf_2 <= _source_stream_conv2d_2_source_25_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_size_buf_3 <= _source_stream_conv2d_2_source_25_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_stride_buf_0 <= _source_stream_conv2d_2_source_25_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_stride_buf_1 <= _source_stream_conv2d_2_source_25_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_stride_buf_2 <= _source_stream_conv2d_2_source_25_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_stride_buf_3 <= _source_stream_conv2d_2_source_25_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_318 <= _stream_conv2d_2_source_25_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_25_idle <= 0;
        _stream_conv2d_2_source_25_source_ram_raddr <= _stream_conv2d_2_source_25_source_pat_all_offset;
        _stream_conv2d_2_source_25_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_0 <= _source_stream_conv2d_2_source_25_pat_cur_offset_0 + _source_stream_conv2d_2_source_25_pat_stride_buf_0;
        _source_stream_conv2d_2_source_25_pat_count_0 <= _source_stream_conv2d_2_source_25_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && (_source_stream_conv2d_2_source_25_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_25_pat_count_0 <= _source_stream_conv2d_2_source_25_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && (_source_stream_conv2d_2_source_25_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_1 <= _source_stream_conv2d_2_source_25_pat_cur_offset_1 + _source_stream_conv2d_2_source_25_pat_stride_buf_1;
        _source_stream_conv2d_2_source_25_pat_count_1 <= _source_stream_conv2d_2_source_25_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && (_source_stream_conv2d_2_source_25_pat_count_0 == 0) && (_source_stream_conv2d_2_source_25_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_25_pat_count_1 <= _source_stream_conv2d_2_source_25_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_2_source_25_pat_count_0 == 0) && (_source_stream_conv2d_2_source_25_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_2 <= _source_stream_conv2d_2_source_25_pat_cur_offset_2 + _source_stream_conv2d_2_source_25_pat_stride_buf_2;
        _source_stream_conv2d_2_source_25_pat_count_2 <= _source_stream_conv2d_2_source_25_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_2_source_25_pat_count_0 == 0) && (_source_stream_conv2d_2_source_25_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_25_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_25_pat_count_2 <= _source_stream_conv2d_2_source_25_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_2_source_25_pat_count_0 == 0) && (_source_stream_conv2d_2_source_25_pat_count_1 == 0) && (_source_stream_conv2d_2_source_25_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_3 <= _source_stream_conv2d_2_source_25_pat_cur_offset_3 + _source_stream_conv2d_2_source_25_pat_stride_buf_3;
        _source_stream_conv2d_2_source_25_pat_count_3 <= _source_stream_conv2d_2_source_25_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_2_source_25_pat_count_0 == 0) && (_source_stream_conv2d_2_source_25_pat_count_1 == 0) && (_source_stream_conv2d_2_source_25_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_25_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_25_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_25_pat_count_3 <= _source_stream_conv2d_2_source_25_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_25_source_ram_renable <= 0;
        _stream_conv2d_2_source_25_idle <= 1;
      end 
      if((_stream_conv2d_2_source_25_source_pat_fsm_5 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_25_source_ram_renable <= 0;
        _stream_conv2d_2_source_25_idle <= 1;
      end 
      if(_set_flag_214) begin
        _stream_conv2d_2_source_26_source_mode <= 5'b10;
        _stream_conv2d_2_source_26_source_offset <= conv2d_2_stream_act_local_6 + conv2d_2_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_214) begin
        _source_stream_conv2d_2_source_26_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_26_pat_stride_0 <= 1;
      end 
      if(_set_flag_214) begin
        _source_stream_conv2d_2_source_26_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_26_pat_stride_1 <= 0;
      end 
      if(_set_flag_214) begin
        _source_stream_conv2d_2_source_26_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_26_pat_stride_2 <= 0;
      end 
      if(_set_flag_214) begin
        _source_stream_conv2d_2_source_26_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_26_pat_stride_3 <= 0;
      end 
      if(_set_flag_214) begin
        _stream_conv2d_2_source_26_source_sel <= 7;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_26_source_offset_buf <= _stream_conv2d_2_source_26_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_count_0 <= _source_stream_conv2d_2_source_26_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_count_1 <= _source_stream_conv2d_2_source_26_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_count_2 <= _source_stream_conv2d_2_source_26_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_count_3 <= _source_stream_conv2d_2_source_26_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_size_buf_0 <= _source_stream_conv2d_2_source_26_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_size_buf_1 <= _source_stream_conv2d_2_source_26_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_size_buf_2 <= _source_stream_conv2d_2_source_26_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_size_buf_3 <= _source_stream_conv2d_2_source_26_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_stride_buf_0 <= _source_stream_conv2d_2_source_26_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_stride_buf_1 <= _source_stream_conv2d_2_source_26_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_stride_buf_2 <= _source_stream_conv2d_2_source_26_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_stride_buf_3 <= _source_stream_conv2d_2_source_26_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_319 <= _stream_conv2d_2_source_26_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_26_idle <= 0;
        _stream_conv2d_2_source_26_source_ram_raddr <= _stream_conv2d_2_source_26_source_pat_all_offset;
        _stream_conv2d_2_source_26_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_0 <= _source_stream_conv2d_2_source_26_pat_cur_offset_0 + _source_stream_conv2d_2_source_26_pat_stride_buf_0;
        _source_stream_conv2d_2_source_26_pat_count_0 <= _source_stream_conv2d_2_source_26_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && (_source_stream_conv2d_2_source_26_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_26_pat_count_0 <= _source_stream_conv2d_2_source_26_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && (_source_stream_conv2d_2_source_26_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_1 <= _source_stream_conv2d_2_source_26_pat_cur_offset_1 + _source_stream_conv2d_2_source_26_pat_stride_buf_1;
        _source_stream_conv2d_2_source_26_pat_count_1 <= _source_stream_conv2d_2_source_26_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && (_source_stream_conv2d_2_source_26_pat_count_0 == 0) && (_source_stream_conv2d_2_source_26_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_26_pat_count_1 <= _source_stream_conv2d_2_source_26_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_2_source_26_pat_count_0 == 0) && (_source_stream_conv2d_2_source_26_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_2 <= _source_stream_conv2d_2_source_26_pat_cur_offset_2 + _source_stream_conv2d_2_source_26_pat_stride_buf_2;
        _source_stream_conv2d_2_source_26_pat_count_2 <= _source_stream_conv2d_2_source_26_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_2_source_26_pat_count_0 == 0) && (_source_stream_conv2d_2_source_26_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_26_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_26_pat_count_2 <= _source_stream_conv2d_2_source_26_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_2_source_26_pat_count_0 == 0) && (_source_stream_conv2d_2_source_26_pat_count_1 == 0) && (_source_stream_conv2d_2_source_26_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_3 <= _source_stream_conv2d_2_source_26_pat_cur_offset_3 + _source_stream_conv2d_2_source_26_pat_stride_buf_3;
        _source_stream_conv2d_2_source_26_pat_count_3 <= _source_stream_conv2d_2_source_26_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_2_source_26_pat_count_0 == 0) && (_source_stream_conv2d_2_source_26_pat_count_1 == 0) && (_source_stream_conv2d_2_source_26_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_26_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_26_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_26_pat_count_3 <= _source_stream_conv2d_2_source_26_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_26_source_ram_renable <= 0;
        _stream_conv2d_2_source_26_idle <= 1;
      end 
      if((_stream_conv2d_2_source_26_source_pat_fsm_6 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_26_source_ram_renable <= 0;
        _stream_conv2d_2_source_26_idle <= 1;
      end 
      if(_set_flag_217) begin
        _stream_conv2d_2_source_27_source_mode <= 5'b10;
        _stream_conv2d_2_source_27_source_offset <= conv2d_2_stream_act_local_7 + conv2d_2_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_217) begin
        _source_stream_conv2d_2_source_27_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_27_pat_stride_0 <= 1;
      end 
      if(_set_flag_217) begin
        _source_stream_conv2d_2_source_27_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_27_pat_stride_1 <= 0;
      end 
      if(_set_flag_217) begin
        _source_stream_conv2d_2_source_27_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_27_pat_stride_2 <= 0;
      end 
      if(_set_flag_217) begin
        _source_stream_conv2d_2_source_27_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_27_pat_stride_3 <= 0;
      end 
      if(_set_flag_217) begin
        _stream_conv2d_2_source_27_source_sel <= 8;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_27_source_offset_buf <= _stream_conv2d_2_source_27_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_count_0 <= _source_stream_conv2d_2_source_27_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_count_1 <= _source_stream_conv2d_2_source_27_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_count_2 <= _source_stream_conv2d_2_source_27_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_count_3 <= _source_stream_conv2d_2_source_27_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_size_buf_0 <= _source_stream_conv2d_2_source_27_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_size_buf_1 <= _source_stream_conv2d_2_source_27_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_size_buf_2 <= _source_stream_conv2d_2_source_27_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_size_buf_3 <= _source_stream_conv2d_2_source_27_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_stride_buf_0 <= _source_stream_conv2d_2_source_27_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_stride_buf_1 <= _source_stream_conv2d_2_source_27_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_stride_buf_2 <= _source_stream_conv2d_2_source_27_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_stride_buf_3 <= _source_stream_conv2d_2_source_27_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_320 <= _stream_conv2d_2_source_27_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_27_idle <= 0;
        _stream_conv2d_2_source_27_source_ram_raddr <= _stream_conv2d_2_source_27_source_pat_all_offset;
        _stream_conv2d_2_source_27_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_0 <= _source_stream_conv2d_2_source_27_pat_cur_offset_0 + _source_stream_conv2d_2_source_27_pat_stride_buf_0;
        _source_stream_conv2d_2_source_27_pat_count_0 <= _source_stream_conv2d_2_source_27_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && (_source_stream_conv2d_2_source_27_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_27_pat_count_0 <= _source_stream_conv2d_2_source_27_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && (_source_stream_conv2d_2_source_27_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_1 <= _source_stream_conv2d_2_source_27_pat_cur_offset_1 + _source_stream_conv2d_2_source_27_pat_stride_buf_1;
        _source_stream_conv2d_2_source_27_pat_count_1 <= _source_stream_conv2d_2_source_27_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && (_source_stream_conv2d_2_source_27_pat_count_0 == 0) && (_source_stream_conv2d_2_source_27_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_27_pat_count_1 <= _source_stream_conv2d_2_source_27_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_2_source_27_pat_count_0 == 0) && (_source_stream_conv2d_2_source_27_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_2 <= _source_stream_conv2d_2_source_27_pat_cur_offset_2 + _source_stream_conv2d_2_source_27_pat_stride_buf_2;
        _source_stream_conv2d_2_source_27_pat_count_2 <= _source_stream_conv2d_2_source_27_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_2_source_27_pat_count_0 == 0) && (_source_stream_conv2d_2_source_27_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_27_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_27_pat_count_2 <= _source_stream_conv2d_2_source_27_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_2_source_27_pat_count_0 == 0) && (_source_stream_conv2d_2_source_27_pat_count_1 == 0) && (_source_stream_conv2d_2_source_27_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_3 <= _source_stream_conv2d_2_source_27_pat_cur_offset_3 + _source_stream_conv2d_2_source_27_pat_stride_buf_3;
        _source_stream_conv2d_2_source_27_pat_count_3 <= _source_stream_conv2d_2_source_27_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_2_source_27_pat_count_0 == 0) && (_source_stream_conv2d_2_source_27_pat_count_1 == 0) && (_source_stream_conv2d_2_source_27_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_27_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_27_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_27_pat_count_3 <= _source_stream_conv2d_2_source_27_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_27_source_ram_renable <= 0;
        _stream_conv2d_2_source_27_idle <= 1;
      end 
      if((_stream_conv2d_2_source_27_source_pat_fsm_7 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_27_source_ram_renable <= 0;
        _stream_conv2d_2_source_27_idle <= 1;
      end 
      if(_set_flag_220) begin
        _stream_conv2d_2_source_28_source_mode <= 5'b10;
        _stream_conv2d_2_source_28_source_offset <= conv2d_2_stream_act_local_8 + conv2d_2_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_220) begin
        _source_stream_conv2d_2_source_28_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_28_pat_stride_0 <= 1;
      end 
      if(_set_flag_220) begin
        _source_stream_conv2d_2_source_28_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_28_pat_stride_1 <= 0;
      end 
      if(_set_flag_220) begin
        _source_stream_conv2d_2_source_28_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_28_pat_stride_2 <= 0;
      end 
      if(_set_flag_220) begin
        _source_stream_conv2d_2_source_28_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_28_pat_stride_3 <= 0;
      end 
      if(_set_flag_220) begin
        _stream_conv2d_2_source_28_source_sel <= 9;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_28_source_offset_buf <= _stream_conv2d_2_source_28_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_count_0 <= _source_stream_conv2d_2_source_28_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_count_1 <= _source_stream_conv2d_2_source_28_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_count_2 <= _source_stream_conv2d_2_source_28_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_count_3 <= _source_stream_conv2d_2_source_28_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_size_buf_0 <= _source_stream_conv2d_2_source_28_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_size_buf_1 <= _source_stream_conv2d_2_source_28_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_size_buf_2 <= _source_stream_conv2d_2_source_28_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_size_buf_3 <= _source_stream_conv2d_2_source_28_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_stride_buf_0 <= _source_stream_conv2d_2_source_28_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_stride_buf_1 <= _source_stream_conv2d_2_source_28_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_stride_buf_2 <= _source_stream_conv2d_2_source_28_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_stride_buf_3 <= _source_stream_conv2d_2_source_28_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_321 <= _stream_conv2d_2_source_28_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_28_idle <= 0;
        _stream_conv2d_2_source_28_source_ram_raddr <= _stream_conv2d_2_source_28_source_pat_all_offset;
        _stream_conv2d_2_source_28_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_0 <= _source_stream_conv2d_2_source_28_pat_cur_offset_0 + _source_stream_conv2d_2_source_28_pat_stride_buf_0;
        _source_stream_conv2d_2_source_28_pat_count_0 <= _source_stream_conv2d_2_source_28_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && (_source_stream_conv2d_2_source_28_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_28_pat_count_0 <= _source_stream_conv2d_2_source_28_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && (_source_stream_conv2d_2_source_28_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_1 <= _source_stream_conv2d_2_source_28_pat_cur_offset_1 + _source_stream_conv2d_2_source_28_pat_stride_buf_1;
        _source_stream_conv2d_2_source_28_pat_count_1 <= _source_stream_conv2d_2_source_28_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && (_source_stream_conv2d_2_source_28_pat_count_0 == 0) && (_source_stream_conv2d_2_source_28_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_28_pat_count_1 <= _source_stream_conv2d_2_source_28_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_2_source_28_pat_count_0 == 0) && (_source_stream_conv2d_2_source_28_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_2 <= _source_stream_conv2d_2_source_28_pat_cur_offset_2 + _source_stream_conv2d_2_source_28_pat_stride_buf_2;
        _source_stream_conv2d_2_source_28_pat_count_2 <= _source_stream_conv2d_2_source_28_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_2_source_28_pat_count_0 == 0) && (_source_stream_conv2d_2_source_28_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_28_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_28_pat_count_2 <= _source_stream_conv2d_2_source_28_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_2_source_28_pat_count_0 == 0) && (_source_stream_conv2d_2_source_28_pat_count_1 == 0) && (_source_stream_conv2d_2_source_28_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_3 <= _source_stream_conv2d_2_source_28_pat_cur_offset_3 + _source_stream_conv2d_2_source_28_pat_stride_buf_3;
        _source_stream_conv2d_2_source_28_pat_count_3 <= _source_stream_conv2d_2_source_28_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_2_source_28_pat_count_0 == 0) && (_source_stream_conv2d_2_source_28_pat_count_1 == 0) && (_source_stream_conv2d_2_source_28_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_28_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_28_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_28_pat_count_3 <= _source_stream_conv2d_2_source_28_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_28_source_ram_renable <= 0;
        _stream_conv2d_2_source_28_idle <= 1;
      end 
      if((_stream_conv2d_2_source_28_source_pat_fsm_8 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_28_source_ram_renable <= 0;
        _stream_conv2d_2_source_28_idle <= 1;
      end 
      if(_set_flag_223) begin
        _stream_conv2d_2_source_29_source_mode <= 5'b10;
        _stream_conv2d_2_source_29_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_223) begin
        _source_stream_conv2d_2_source_29_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_29_pat_stride_0 <= 1;
      end 
      if(_set_flag_223) begin
        _source_stream_conv2d_2_source_29_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_29_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_223) begin
        _source_stream_conv2d_2_source_29_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_29_pat_stride_2 <= 0;
      end 
      if(_set_flag_223) begin
        _source_stream_conv2d_2_source_29_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_29_pat_stride_3 <= 0;
      end 
      if(_set_flag_223) begin
        _stream_conv2d_2_source_29_source_sel <= 10;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_29_source_offset_buf <= _stream_conv2d_2_source_29_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_count_0 <= _source_stream_conv2d_2_source_29_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_count_1 <= _source_stream_conv2d_2_source_29_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_count_2 <= _source_stream_conv2d_2_source_29_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_count_3 <= _source_stream_conv2d_2_source_29_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_size_buf_0 <= _source_stream_conv2d_2_source_29_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_size_buf_1 <= _source_stream_conv2d_2_source_29_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_size_buf_2 <= _source_stream_conv2d_2_source_29_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_size_buf_3 <= _source_stream_conv2d_2_source_29_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_stride_buf_0 <= _source_stream_conv2d_2_source_29_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_stride_buf_1 <= _source_stream_conv2d_2_source_29_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_stride_buf_2 <= _source_stream_conv2d_2_source_29_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_stride_buf_3 <= _source_stream_conv2d_2_source_29_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_547 <= _stream_conv2d_2_source_29_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_29_idle <= 0;
        _stream_conv2d_2_source_29_source_ram_raddr <= _stream_conv2d_2_source_29_source_pat_all_offset;
        _stream_conv2d_2_source_29_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_0 <= _source_stream_conv2d_2_source_29_pat_cur_offset_0 + _source_stream_conv2d_2_source_29_pat_stride_buf_0;
        _source_stream_conv2d_2_source_29_pat_count_0 <= _source_stream_conv2d_2_source_29_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && (_source_stream_conv2d_2_source_29_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_29_pat_count_0 <= _source_stream_conv2d_2_source_29_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && (_source_stream_conv2d_2_source_29_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_1 <= _source_stream_conv2d_2_source_29_pat_cur_offset_1 + _source_stream_conv2d_2_source_29_pat_stride_buf_1;
        _source_stream_conv2d_2_source_29_pat_count_1 <= _source_stream_conv2d_2_source_29_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && (_source_stream_conv2d_2_source_29_pat_count_0 == 0) && (_source_stream_conv2d_2_source_29_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_29_pat_count_1 <= _source_stream_conv2d_2_source_29_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_2_source_29_pat_count_0 == 0) && (_source_stream_conv2d_2_source_29_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_2 <= _source_stream_conv2d_2_source_29_pat_cur_offset_2 + _source_stream_conv2d_2_source_29_pat_stride_buf_2;
        _source_stream_conv2d_2_source_29_pat_count_2 <= _source_stream_conv2d_2_source_29_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_2_source_29_pat_count_0 == 0) && (_source_stream_conv2d_2_source_29_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_29_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_29_pat_count_2 <= _source_stream_conv2d_2_source_29_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_2_source_29_pat_count_0 == 0) && (_source_stream_conv2d_2_source_29_pat_count_1 == 0) && (_source_stream_conv2d_2_source_29_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_3 <= _source_stream_conv2d_2_source_29_pat_cur_offset_3 + _source_stream_conv2d_2_source_29_pat_stride_buf_3;
        _source_stream_conv2d_2_source_29_pat_count_3 <= _source_stream_conv2d_2_source_29_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_2_source_29_pat_count_0 == 0) && (_source_stream_conv2d_2_source_29_pat_count_1 == 0) && (_source_stream_conv2d_2_source_29_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_29_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_29_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_29_pat_count_3 <= _source_stream_conv2d_2_source_29_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_29_source_ram_renable <= 0;
        _stream_conv2d_2_source_29_idle <= 1;
      end 
      if((_stream_conv2d_2_source_29_source_pat_fsm_9 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_29_source_ram_renable <= 0;
        _stream_conv2d_2_source_29_idle <= 1;
      end 
      if(_set_flag_226) begin
        _stream_conv2d_2_source_30_source_mode <= 5'b10;
        _stream_conv2d_2_source_30_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_226) begin
        _source_stream_conv2d_2_source_30_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_30_pat_stride_0 <= 1;
      end 
      if(_set_flag_226) begin
        _source_stream_conv2d_2_source_30_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_30_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_226) begin
        _source_stream_conv2d_2_source_30_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_30_pat_stride_2 <= 0;
      end 
      if(_set_flag_226) begin
        _source_stream_conv2d_2_source_30_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_30_pat_stride_3 <= 0;
      end 
      if(_set_flag_226) begin
        _stream_conv2d_2_source_30_source_sel <= 11;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_30_source_offset_buf <= _stream_conv2d_2_source_30_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_count_0 <= _source_stream_conv2d_2_source_30_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_count_1 <= _source_stream_conv2d_2_source_30_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_count_2 <= _source_stream_conv2d_2_source_30_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_count_3 <= _source_stream_conv2d_2_source_30_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_size_buf_0 <= _source_stream_conv2d_2_source_30_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_size_buf_1 <= _source_stream_conv2d_2_source_30_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_size_buf_2 <= _source_stream_conv2d_2_source_30_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_size_buf_3 <= _source_stream_conv2d_2_source_30_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_stride_buf_0 <= _source_stream_conv2d_2_source_30_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_stride_buf_1 <= _source_stream_conv2d_2_source_30_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_stride_buf_2 <= _source_stream_conv2d_2_source_30_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_stride_buf_3 <= _source_stream_conv2d_2_source_30_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_548 <= _stream_conv2d_2_source_30_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_30_idle <= 0;
        _stream_conv2d_2_source_30_source_ram_raddr <= _stream_conv2d_2_source_30_source_pat_all_offset;
        _stream_conv2d_2_source_30_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_0 <= _source_stream_conv2d_2_source_30_pat_cur_offset_0 + _source_stream_conv2d_2_source_30_pat_stride_buf_0;
        _source_stream_conv2d_2_source_30_pat_count_0 <= _source_stream_conv2d_2_source_30_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && (_source_stream_conv2d_2_source_30_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_30_pat_count_0 <= _source_stream_conv2d_2_source_30_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && (_source_stream_conv2d_2_source_30_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_1 <= _source_stream_conv2d_2_source_30_pat_cur_offset_1 + _source_stream_conv2d_2_source_30_pat_stride_buf_1;
        _source_stream_conv2d_2_source_30_pat_count_1 <= _source_stream_conv2d_2_source_30_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && (_source_stream_conv2d_2_source_30_pat_count_0 == 0) && (_source_stream_conv2d_2_source_30_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_30_pat_count_1 <= _source_stream_conv2d_2_source_30_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_2_source_30_pat_count_0 == 0) && (_source_stream_conv2d_2_source_30_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_2 <= _source_stream_conv2d_2_source_30_pat_cur_offset_2 + _source_stream_conv2d_2_source_30_pat_stride_buf_2;
        _source_stream_conv2d_2_source_30_pat_count_2 <= _source_stream_conv2d_2_source_30_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_2_source_30_pat_count_0 == 0) && (_source_stream_conv2d_2_source_30_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_30_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_30_pat_count_2 <= _source_stream_conv2d_2_source_30_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_2_source_30_pat_count_0 == 0) && (_source_stream_conv2d_2_source_30_pat_count_1 == 0) && (_source_stream_conv2d_2_source_30_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_3 <= _source_stream_conv2d_2_source_30_pat_cur_offset_3 + _source_stream_conv2d_2_source_30_pat_stride_buf_3;
        _source_stream_conv2d_2_source_30_pat_count_3 <= _source_stream_conv2d_2_source_30_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_2_source_30_pat_count_0 == 0) && (_source_stream_conv2d_2_source_30_pat_count_1 == 0) && (_source_stream_conv2d_2_source_30_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_30_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_30_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_30_pat_count_3 <= _source_stream_conv2d_2_source_30_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_30_source_ram_renable <= 0;
        _stream_conv2d_2_source_30_idle <= 1;
      end 
      if((_stream_conv2d_2_source_30_source_pat_fsm_10 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_30_source_ram_renable <= 0;
        _stream_conv2d_2_source_30_idle <= 1;
      end 
      if(_set_flag_229) begin
        _stream_conv2d_2_source_31_source_mode <= 5'b10;
        _stream_conv2d_2_source_31_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_229) begin
        _source_stream_conv2d_2_source_31_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_31_pat_stride_0 <= 1;
      end 
      if(_set_flag_229) begin
        _source_stream_conv2d_2_source_31_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_31_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_229) begin
        _source_stream_conv2d_2_source_31_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_31_pat_stride_2 <= 0;
      end 
      if(_set_flag_229) begin
        _source_stream_conv2d_2_source_31_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_31_pat_stride_3 <= 0;
      end 
      if(_set_flag_229) begin
        _stream_conv2d_2_source_31_source_sel <= 12;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_31_source_offset_buf <= _stream_conv2d_2_source_31_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_count_0 <= _source_stream_conv2d_2_source_31_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_count_1 <= _source_stream_conv2d_2_source_31_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_count_2 <= _source_stream_conv2d_2_source_31_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_count_3 <= _source_stream_conv2d_2_source_31_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_size_buf_0 <= _source_stream_conv2d_2_source_31_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_size_buf_1 <= _source_stream_conv2d_2_source_31_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_size_buf_2 <= _source_stream_conv2d_2_source_31_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_size_buf_3 <= _source_stream_conv2d_2_source_31_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_stride_buf_0 <= _source_stream_conv2d_2_source_31_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_stride_buf_1 <= _source_stream_conv2d_2_source_31_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_stride_buf_2 <= _source_stream_conv2d_2_source_31_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_stride_buf_3 <= _source_stream_conv2d_2_source_31_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_549 <= _stream_conv2d_2_source_31_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_31_idle <= 0;
        _stream_conv2d_2_source_31_source_ram_raddr <= _stream_conv2d_2_source_31_source_pat_all_offset;
        _stream_conv2d_2_source_31_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_0 <= _source_stream_conv2d_2_source_31_pat_cur_offset_0 + _source_stream_conv2d_2_source_31_pat_stride_buf_0;
        _source_stream_conv2d_2_source_31_pat_count_0 <= _source_stream_conv2d_2_source_31_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && (_source_stream_conv2d_2_source_31_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_31_pat_count_0 <= _source_stream_conv2d_2_source_31_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && (_source_stream_conv2d_2_source_31_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_1 <= _source_stream_conv2d_2_source_31_pat_cur_offset_1 + _source_stream_conv2d_2_source_31_pat_stride_buf_1;
        _source_stream_conv2d_2_source_31_pat_count_1 <= _source_stream_conv2d_2_source_31_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && (_source_stream_conv2d_2_source_31_pat_count_0 == 0) && (_source_stream_conv2d_2_source_31_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_31_pat_count_1 <= _source_stream_conv2d_2_source_31_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_2_source_31_pat_count_0 == 0) && (_source_stream_conv2d_2_source_31_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_2 <= _source_stream_conv2d_2_source_31_pat_cur_offset_2 + _source_stream_conv2d_2_source_31_pat_stride_buf_2;
        _source_stream_conv2d_2_source_31_pat_count_2 <= _source_stream_conv2d_2_source_31_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_2_source_31_pat_count_0 == 0) && (_source_stream_conv2d_2_source_31_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_31_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_31_pat_count_2 <= _source_stream_conv2d_2_source_31_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_2_source_31_pat_count_0 == 0) && (_source_stream_conv2d_2_source_31_pat_count_1 == 0) && (_source_stream_conv2d_2_source_31_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_3 <= _source_stream_conv2d_2_source_31_pat_cur_offset_3 + _source_stream_conv2d_2_source_31_pat_stride_buf_3;
        _source_stream_conv2d_2_source_31_pat_count_3 <= _source_stream_conv2d_2_source_31_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_2_source_31_pat_count_0 == 0) && (_source_stream_conv2d_2_source_31_pat_count_1 == 0) && (_source_stream_conv2d_2_source_31_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_31_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_31_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_31_pat_count_3 <= _source_stream_conv2d_2_source_31_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_31_source_ram_renable <= 0;
        _stream_conv2d_2_source_31_idle <= 1;
      end 
      if((_stream_conv2d_2_source_31_source_pat_fsm_11 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_31_source_ram_renable <= 0;
        _stream_conv2d_2_source_31_idle <= 1;
      end 
      if(_set_flag_232) begin
        _stream_conv2d_2_source_32_source_mode <= 5'b10;
        _stream_conv2d_2_source_32_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_232) begin
        _source_stream_conv2d_2_source_32_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_32_pat_stride_0 <= 1;
      end 
      if(_set_flag_232) begin
        _source_stream_conv2d_2_source_32_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_32_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_232) begin
        _source_stream_conv2d_2_source_32_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_32_pat_stride_2 <= 0;
      end 
      if(_set_flag_232) begin
        _source_stream_conv2d_2_source_32_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_32_pat_stride_3 <= 0;
      end 
      if(_set_flag_232) begin
        _stream_conv2d_2_source_32_source_sel <= 13;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_32_source_offset_buf <= _stream_conv2d_2_source_32_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_count_0 <= _source_stream_conv2d_2_source_32_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_count_1 <= _source_stream_conv2d_2_source_32_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_count_2 <= _source_stream_conv2d_2_source_32_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_count_3 <= _source_stream_conv2d_2_source_32_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_size_buf_0 <= _source_stream_conv2d_2_source_32_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_size_buf_1 <= _source_stream_conv2d_2_source_32_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_size_buf_2 <= _source_stream_conv2d_2_source_32_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_size_buf_3 <= _source_stream_conv2d_2_source_32_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_stride_buf_0 <= _source_stream_conv2d_2_source_32_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_stride_buf_1 <= _source_stream_conv2d_2_source_32_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_stride_buf_2 <= _source_stream_conv2d_2_source_32_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_stride_buf_3 <= _source_stream_conv2d_2_source_32_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_550 <= _stream_conv2d_2_source_32_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_32_idle <= 0;
        _stream_conv2d_2_source_32_source_ram_raddr <= _stream_conv2d_2_source_32_source_pat_all_offset;
        _stream_conv2d_2_source_32_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_0 <= _source_stream_conv2d_2_source_32_pat_cur_offset_0 + _source_stream_conv2d_2_source_32_pat_stride_buf_0;
        _source_stream_conv2d_2_source_32_pat_count_0 <= _source_stream_conv2d_2_source_32_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && (_source_stream_conv2d_2_source_32_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_32_pat_count_0 <= _source_stream_conv2d_2_source_32_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && (_source_stream_conv2d_2_source_32_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_1 <= _source_stream_conv2d_2_source_32_pat_cur_offset_1 + _source_stream_conv2d_2_source_32_pat_stride_buf_1;
        _source_stream_conv2d_2_source_32_pat_count_1 <= _source_stream_conv2d_2_source_32_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && (_source_stream_conv2d_2_source_32_pat_count_0 == 0) && (_source_stream_conv2d_2_source_32_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_32_pat_count_1 <= _source_stream_conv2d_2_source_32_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_2_source_32_pat_count_0 == 0) && (_source_stream_conv2d_2_source_32_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_2 <= _source_stream_conv2d_2_source_32_pat_cur_offset_2 + _source_stream_conv2d_2_source_32_pat_stride_buf_2;
        _source_stream_conv2d_2_source_32_pat_count_2 <= _source_stream_conv2d_2_source_32_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_2_source_32_pat_count_0 == 0) && (_source_stream_conv2d_2_source_32_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_32_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_32_pat_count_2 <= _source_stream_conv2d_2_source_32_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_2_source_32_pat_count_0 == 0) && (_source_stream_conv2d_2_source_32_pat_count_1 == 0) && (_source_stream_conv2d_2_source_32_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_3 <= _source_stream_conv2d_2_source_32_pat_cur_offset_3 + _source_stream_conv2d_2_source_32_pat_stride_buf_3;
        _source_stream_conv2d_2_source_32_pat_count_3 <= _source_stream_conv2d_2_source_32_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_2_source_32_pat_count_0 == 0) && (_source_stream_conv2d_2_source_32_pat_count_1 == 0) && (_source_stream_conv2d_2_source_32_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_32_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_32_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_32_pat_count_3 <= _source_stream_conv2d_2_source_32_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_32_source_ram_renable <= 0;
        _stream_conv2d_2_source_32_idle <= 1;
      end 
      if((_stream_conv2d_2_source_32_source_pat_fsm_12 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_32_source_ram_renable <= 0;
        _stream_conv2d_2_source_32_idle <= 1;
      end 
      if(_set_flag_235) begin
        _stream_conv2d_2_source_33_source_mode <= 5'b10;
        _stream_conv2d_2_source_33_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_235) begin
        _source_stream_conv2d_2_source_33_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_33_pat_stride_0 <= 1;
      end 
      if(_set_flag_235) begin
        _source_stream_conv2d_2_source_33_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_33_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_235) begin
        _source_stream_conv2d_2_source_33_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_33_pat_stride_2 <= 0;
      end 
      if(_set_flag_235) begin
        _source_stream_conv2d_2_source_33_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_33_pat_stride_3 <= 0;
      end 
      if(_set_flag_235) begin
        _stream_conv2d_2_source_33_source_sel <= 14;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_33_source_offset_buf <= _stream_conv2d_2_source_33_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_count_0 <= _source_stream_conv2d_2_source_33_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_count_1 <= _source_stream_conv2d_2_source_33_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_count_2 <= _source_stream_conv2d_2_source_33_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_count_3 <= _source_stream_conv2d_2_source_33_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_size_buf_0 <= _source_stream_conv2d_2_source_33_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_size_buf_1 <= _source_stream_conv2d_2_source_33_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_size_buf_2 <= _source_stream_conv2d_2_source_33_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_size_buf_3 <= _source_stream_conv2d_2_source_33_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_stride_buf_0 <= _source_stream_conv2d_2_source_33_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_stride_buf_1 <= _source_stream_conv2d_2_source_33_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_stride_buf_2 <= _source_stream_conv2d_2_source_33_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_stride_buf_3 <= _source_stream_conv2d_2_source_33_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_551 <= _stream_conv2d_2_source_33_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_33_idle <= 0;
        _stream_conv2d_2_source_33_source_ram_raddr <= _stream_conv2d_2_source_33_source_pat_all_offset;
        _stream_conv2d_2_source_33_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_0 <= _source_stream_conv2d_2_source_33_pat_cur_offset_0 + _source_stream_conv2d_2_source_33_pat_stride_buf_0;
        _source_stream_conv2d_2_source_33_pat_count_0 <= _source_stream_conv2d_2_source_33_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && (_source_stream_conv2d_2_source_33_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_33_pat_count_0 <= _source_stream_conv2d_2_source_33_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && (_source_stream_conv2d_2_source_33_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_1 <= _source_stream_conv2d_2_source_33_pat_cur_offset_1 + _source_stream_conv2d_2_source_33_pat_stride_buf_1;
        _source_stream_conv2d_2_source_33_pat_count_1 <= _source_stream_conv2d_2_source_33_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && (_source_stream_conv2d_2_source_33_pat_count_0 == 0) && (_source_stream_conv2d_2_source_33_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_33_pat_count_1 <= _source_stream_conv2d_2_source_33_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_2_source_33_pat_count_0 == 0) && (_source_stream_conv2d_2_source_33_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_2 <= _source_stream_conv2d_2_source_33_pat_cur_offset_2 + _source_stream_conv2d_2_source_33_pat_stride_buf_2;
        _source_stream_conv2d_2_source_33_pat_count_2 <= _source_stream_conv2d_2_source_33_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_2_source_33_pat_count_0 == 0) && (_source_stream_conv2d_2_source_33_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_33_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_33_pat_count_2 <= _source_stream_conv2d_2_source_33_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_2_source_33_pat_count_0 == 0) && (_source_stream_conv2d_2_source_33_pat_count_1 == 0) && (_source_stream_conv2d_2_source_33_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_3 <= _source_stream_conv2d_2_source_33_pat_cur_offset_3 + _source_stream_conv2d_2_source_33_pat_stride_buf_3;
        _source_stream_conv2d_2_source_33_pat_count_3 <= _source_stream_conv2d_2_source_33_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_2_source_33_pat_count_0 == 0) && (_source_stream_conv2d_2_source_33_pat_count_1 == 0) && (_source_stream_conv2d_2_source_33_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_33_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_33_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_33_pat_count_3 <= _source_stream_conv2d_2_source_33_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_33_source_ram_renable <= 0;
        _stream_conv2d_2_source_33_idle <= 1;
      end 
      if((_stream_conv2d_2_source_33_source_pat_fsm_13 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_33_source_ram_renable <= 0;
        _stream_conv2d_2_source_33_idle <= 1;
      end 
      if(_set_flag_238) begin
        _stream_conv2d_2_source_34_source_mode <= 5'b10;
        _stream_conv2d_2_source_34_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_238) begin
        _source_stream_conv2d_2_source_34_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_34_pat_stride_0 <= 1;
      end 
      if(_set_flag_238) begin
        _source_stream_conv2d_2_source_34_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_34_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_238) begin
        _source_stream_conv2d_2_source_34_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_34_pat_stride_2 <= 0;
      end 
      if(_set_flag_238) begin
        _source_stream_conv2d_2_source_34_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_34_pat_stride_3 <= 0;
      end 
      if(_set_flag_238) begin
        _stream_conv2d_2_source_34_source_sel <= 15;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_34_source_offset_buf <= _stream_conv2d_2_source_34_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_count_0 <= _source_stream_conv2d_2_source_34_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_count_1 <= _source_stream_conv2d_2_source_34_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_count_2 <= _source_stream_conv2d_2_source_34_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_count_3 <= _source_stream_conv2d_2_source_34_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_size_buf_0 <= _source_stream_conv2d_2_source_34_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_size_buf_1 <= _source_stream_conv2d_2_source_34_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_size_buf_2 <= _source_stream_conv2d_2_source_34_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_size_buf_3 <= _source_stream_conv2d_2_source_34_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_stride_buf_0 <= _source_stream_conv2d_2_source_34_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_stride_buf_1 <= _source_stream_conv2d_2_source_34_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_stride_buf_2 <= _source_stream_conv2d_2_source_34_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_stride_buf_3 <= _source_stream_conv2d_2_source_34_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_552 <= _stream_conv2d_2_source_34_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_34_idle <= 0;
        _stream_conv2d_2_source_34_source_ram_raddr <= _stream_conv2d_2_source_34_source_pat_all_offset;
        _stream_conv2d_2_source_34_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_0 <= _source_stream_conv2d_2_source_34_pat_cur_offset_0 + _source_stream_conv2d_2_source_34_pat_stride_buf_0;
        _source_stream_conv2d_2_source_34_pat_count_0 <= _source_stream_conv2d_2_source_34_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && (_source_stream_conv2d_2_source_34_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_34_pat_count_0 <= _source_stream_conv2d_2_source_34_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && (_source_stream_conv2d_2_source_34_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_1 <= _source_stream_conv2d_2_source_34_pat_cur_offset_1 + _source_stream_conv2d_2_source_34_pat_stride_buf_1;
        _source_stream_conv2d_2_source_34_pat_count_1 <= _source_stream_conv2d_2_source_34_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && (_source_stream_conv2d_2_source_34_pat_count_0 == 0) && (_source_stream_conv2d_2_source_34_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_34_pat_count_1 <= _source_stream_conv2d_2_source_34_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_2_source_34_pat_count_0 == 0) && (_source_stream_conv2d_2_source_34_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_2 <= _source_stream_conv2d_2_source_34_pat_cur_offset_2 + _source_stream_conv2d_2_source_34_pat_stride_buf_2;
        _source_stream_conv2d_2_source_34_pat_count_2 <= _source_stream_conv2d_2_source_34_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_2_source_34_pat_count_0 == 0) && (_source_stream_conv2d_2_source_34_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_34_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_34_pat_count_2 <= _source_stream_conv2d_2_source_34_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_2_source_34_pat_count_0 == 0) && (_source_stream_conv2d_2_source_34_pat_count_1 == 0) && (_source_stream_conv2d_2_source_34_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_3 <= _source_stream_conv2d_2_source_34_pat_cur_offset_3 + _source_stream_conv2d_2_source_34_pat_stride_buf_3;
        _source_stream_conv2d_2_source_34_pat_count_3 <= _source_stream_conv2d_2_source_34_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_2_source_34_pat_count_0 == 0) && (_source_stream_conv2d_2_source_34_pat_count_1 == 0) && (_source_stream_conv2d_2_source_34_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_34_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_34_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_34_pat_count_3 <= _source_stream_conv2d_2_source_34_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_34_source_ram_renable <= 0;
        _stream_conv2d_2_source_34_idle <= 1;
      end 
      if((_stream_conv2d_2_source_34_source_pat_fsm_14 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_34_source_ram_renable <= 0;
        _stream_conv2d_2_source_34_idle <= 1;
      end 
      if(_set_flag_241) begin
        _stream_conv2d_2_source_35_source_mode <= 5'b10;
        _stream_conv2d_2_source_35_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_2_source_35_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_35_pat_stride_0 <= 1;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_2_source_35_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_35_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_2_source_35_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_35_pat_stride_2 <= 0;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_2_source_35_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_35_pat_stride_3 <= 0;
      end 
      if(_set_flag_241) begin
        _stream_conv2d_2_source_35_source_sel <= 16;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_35_source_offset_buf <= _stream_conv2d_2_source_35_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_count_0 <= _source_stream_conv2d_2_source_35_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_count_1 <= _source_stream_conv2d_2_source_35_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_count_2 <= _source_stream_conv2d_2_source_35_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_count_3 <= _source_stream_conv2d_2_source_35_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_size_buf_0 <= _source_stream_conv2d_2_source_35_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_size_buf_1 <= _source_stream_conv2d_2_source_35_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_size_buf_2 <= _source_stream_conv2d_2_source_35_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_size_buf_3 <= _source_stream_conv2d_2_source_35_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_stride_buf_0 <= _source_stream_conv2d_2_source_35_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_stride_buf_1 <= _source_stream_conv2d_2_source_35_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_stride_buf_2 <= _source_stream_conv2d_2_source_35_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_stride_buf_3 <= _source_stream_conv2d_2_source_35_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_553 <= _stream_conv2d_2_source_35_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_35_idle <= 0;
        _stream_conv2d_2_source_35_source_ram_raddr <= _stream_conv2d_2_source_35_source_pat_all_offset;
        _stream_conv2d_2_source_35_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_0 <= _source_stream_conv2d_2_source_35_pat_cur_offset_0 + _source_stream_conv2d_2_source_35_pat_stride_buf_0;
        _source_stream_conv2d_2_source_35_pat_count_0 <= _source_stream_conv2d_2_source_35_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && (_source_stream_conv2d_2_source_35_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_35_pat_count_0 <= _source_stream_conv2d_2_source_35_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && (_source_stream_conv2d_2_source_35_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_1 <= _source_stream_conv2d_2_source_35_pat_cur_offset_1 + _source_stream_conv2d_2_source_35_pat_stride_buf_1;
        _source_stream_conv2d_2_source_35_pat_count_1 <= _source_stream_conv2d_2_source_35_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && (_source_stream_conv2d_2_source_35_pat_count_0 == 0) && (_source_stream_conv2d_2_source_35_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_35_pat_count_1 <= _source_stream_conv2d_2_source_35_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_2_source_35_pat_count_0 == 0) && (_source_stream_conv2d_2_source_35_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_2 <= _source_stream_conv2d_2_source_35_pat_cur_offset_2 + _source_stream_conv2d_2_source_35_pat_stride_buf_2;
        _source_stream_conv2d_2_source_35_pat_count_2 <= _source_stream_conv2d_2_source_35_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_2_source_35_pat_count_0 == 0) && (_source_stream_conv2d_2_source_35_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_35_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_35_pat_count_2 <= _source_stream_conv2d_2_source_35_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_2_source_35_pat_count_0 == 0) && (_source_stream_conv2d_2_source_35_pat_count_1 == 0) && (_source_stream_conv2d_2_source_35_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_3 <= _source_stream_conv2d_2_source_35_pat_cur_offset_3 + _source_stream_conv2d_2_source_35_pat_stride_buf_3;
        _source_stream_conv2d_2_source_35_pat_count_3 <= _source_stream_conv2d_2_source_35_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_2_source_35_pat_count_0 == 0) && (_source_stream_conv2d_2_source_35_pat_count_1 == 0) && (_source_stream_conv2d_2_source_35_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_35_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_35_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_35_pat_count_3 <= _source_stream_conv2d_2_source_35_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_35_source_ram_renable <= 0;
        _stream_conv2d_2_source_35_idle <= 1;
      end 
      if((_stream_conv2d_2_source_35_source_pat_fsm_15 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_35_source_ram_renable <= 0;
        _stream_conv2d_2_source_35_idle <= 1;
      end 
      if(_set_flag_244) begin
        _stream_conv2d_2_source_36_source_mode <= 5'b10;
        _stream_conv2d_2_source_36_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_2_source_36_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_36_pat_stride_0 <= 1;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_2_source_36_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_36_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_2_source_36_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_36_pat_stride_2 <= 0;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_2_source_36_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_36_pat_stride_3 <= 0;
      end 
      if(_set_flag_244) begin
        _stream_conv2d_2_source_36_source_sel <= 17;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_36_source_offset_buf <= _stream_conv2d_2_source_36_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_count_0 <= _source_stream_conv2d_2_source_36_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_count_1 <= _source_stream_conv2d_2_source_36_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_count_2 <= _source_stream_conv2d_2_source_36_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_count_3 <= _source_stream_conv2d_2_source_36_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_size_buf_0 <= _source_stream_conv2d_2_source_36_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_size_buf_1 <= _source_stream_conv2d_2_source_36_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_size_buf_2 <= _source_stream_conv2d_2_source_36_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_size_buf_3 <= _source_stream_conv2d_2_source_36_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_stride_buf_0 <= _source_stream_conv2d_2_source_36_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_stride_buf_1 <= _source_stream_conv2d_2_source_36_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_stride_buf_2 <= _source_stream_conv2d_2_source_36_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_stride_buf_3 <= _source_stream_conv2d_2_source_36_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_554 <= _stream_conv2d_2_source_36_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_36_idle <= 0;
        _stream_conv2d_2_source_36_source_ram_raddr <= _stream_conv2d_2_source_36_source_pat_all_offset;
        _stream_conv2d_2_source_36_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_0 <= _source_stream_conv2d_2_source_36_pat_cur_offset_0 + _source_stream_conv2d_2_source_36_pat_stride_buf_0;
        _source_stream_conv2d_2_source_36_pat_count_0 <= _source_stream_conv2d_2_source_36_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && (_source_stream_conv2d_2_source_36_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_36_pat_count_0 <= _source_stream_conv2d_2_source_36_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && (_source_stream_conv2d_2_source_36_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_1 <= _source_stream_conv2d_2_source_36_pat_cur_offset_1 + _source_stream_conv2d_2_source_36_pat_stride_buf_1;
        _source_stream_conv2d_2_source_36_pat_count_1 <= _source_stream_conv2d_2_source_36_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && (_source_stream_conv2d_2_source_36_pat_count_0 == 0) && (_source_stream_conv2d_2_source_36_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_36_pat_count_1 <= _source_stream_conv2d_2_source_36_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_2_source_36_pat_count_0 == 0) && (_source_stream_conv2d_2_source_36_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_2 <= _source_stream_conv2d_2_source_36_pat_cur_offset_2 + _source_stream_conv2d_2_source_36_pat_stride_buf_2;
        _source_stream_conv2d_2_source_36_pat_count_2 <= _source_stream_conv2d_2_source_36_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_2_source_36_pat_count_0 == 0) && (_source_stream_conv2d_2_source_36_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_36_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_36_pat_count_2 <= _source_stream_conv2d_2_source_36_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_2_source_36_pat_count_0 == 0) && (_source_stream_conv2d_2_source_36_pat_count_1 == 0) && (_source_stream_conv2d_2_source_36_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_3 <= _source_stream_conv2d_2_source_36_pat_cur_offset_3 + _source_stream_conv2d_2_source_36_pat_stride_buf_3;
        _source_stream_conv2d_2_source_36_pat_count_3 <= _source_stream_conv2d_2_source_36_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_2_source_36_pat_count_0 == 0) && (_source_stream_conv2d_2_source_36_pat_count_1 == 0) && (_source_stream_conv2d_2_source_36_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_36_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_36_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_36_pat_count_3 <= _source_stream_conv2d_2_source_36_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_36_source_ram_renable <= 0;
        _stream_conv2d_2_source_36_idle <= 1;
      end 
      if((_stream_conv2d_2_source_36_source_pat_fsm_16 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_36_source_ram_renable <= 0;
        _stream_conv2d_2_source_36_idle <= 1;
      end 
      if(_set_flag_247) begin
        _stream_conv2d_2_source_37_source_mode <= 5'b10;
        _stream_conv2d_2_source_37_source_offset <= conv2d_2_filter_page_comp_offset_buf;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_2_source_37_pat_size_0 <= cparam_conv2d_2_stream_reduce_size;
        _source_stream_conv2d_2_source_37_pat_stride_0 <= 1;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_2_source_37_pat_size_1 <= conv2d_2_next_stream_num_ops;
        _source_stream_conv2d_2_source_37_pat_stride_1 <= cparam_conv2d_2_stream_aligned_reduce_size;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_2_source_37_pat_size_2 <= 1;
        _source_stream_conv2d_2_source_37_pat_stride_2 <= 0;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_2_source_37_pat_size_3 <= 1;
        _source_stream_conv2d_2_source_37_pat_stride_3 <= 0;
      end 
      if(_set_flag_247) begin
        _stream_conv2d_2_source_37_source_sel <= 18;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_37_source_offset_buf <= _stream_conv2d_2_source_37_source_offset;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_count_0 <= _source_stream_conv2d_2_source_37_pat_size_0 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_count_1 <= _source_stream_conv2d_2_source_37_pat_size_1 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_count_2 <= _source_stream_conv2d_2_source_37_pat_size_2 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_count_3 <= _source_stream_conv2d_2_source_37_pat_size_3 - 1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_size_buf_0 <= _source_stream_conv2d_2_source_37_pat_size_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_size_buf_1 <= _source_stream_conv2d_2_source_37_pat_size_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_size_buf_2 <= _source_stream_conv2d_2_source_37_pat_size_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_size_buf_3 <= _source_stream_conv2d_2_source_37_pat_size_3;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_stride_buf_0 <= _source_stream_conv2d_2_source_37_pat_stride_0;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_stride_buf_1 <= _source_stream_conv2d_2_source_37_pat_stride_1;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_stride_buf_2 <= _source_stream_conv2d_2_source_37_pat_stride_2;
      end 
      if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_stride_buf_3 <= _source_stream_conv2d_2_source_37_pat_stride_3;
      end 
      if(_stream_conv2d_2_stream_oready && _stream_conv2d_2_source_busy && _stream_conv2d_2_is_root) begin
        __variable_wdata_555 <= _stream_conv2d_2_source_37_source_ram_rdata;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_37_idle <= 0;
        _stream_conv2d_2_source_37_source_ram_raddr <= _stream_conv2d_2_source_37_source_pat_all_offset;
        _stream_conv2d_2_source_37_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_0 <= _source_stream_conv2d_2_source_37_pat_cur_offset_0 + _source_stream_conv2d_2_source_37_pat_stride_buf_0;
        _source_stream_conv2d_2_source_37_pat_count_0 <= _source_stream_conv2d_2_source_37_pat_count_0 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && (_source_stream_conv2d_2_source_37_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_2_source_37_pat_count_0 <= _source_stream_conv2d_2_source_37_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && (_source_stream_conv2d_2_source_37_pat_count_0 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_1 <= _source_stream_conv2d_2_source_37_pat_cur_offset_1 + _source_stream_conv2d_2_source_37_pat_stride_buf_1;
        _source_stream_conv2d_2_source_37_pat_count_1 <= _source_stream_conv2d_2_source_37_pat_count_1 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && (_source_stream_conv2d_2_source_37_pat_count_0 == 0) && (_source_stream_conv2d_2_source_37_pat_count_1 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_2_source_37_pat_count_1 <= _source_stream_conv2d_2_source_37_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_2_source_37_pat_count_0 == 0) && (_source_stream_conv2d_2_source_37_pat_count_1 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_2 <= _source_stream_conv2d_2_source_37_pat_cur_offset_2 + _source_stream_conv2d_2_source_37_pat_stride_buf_2;
        _source_stream_conv2d_2_source_37_pat_count_2 <= _source_stream_conv2d_2_source_37_pat_count_2 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_2_source_37_pat_count_0 == 0) && (_source_stream_conv2d_2_source_37_pat_count_1 == 0)) && (_source_stream_conv2d_2_source_37_pat_count_2 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_2_source_37_pat_count_2 <= _source_stream_conv2d_2_source_37_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_2_source_37_pat_count_0 == 0) && (_source_stream_conv2d_2_source_37_pat_count_1 == 0) && (_source_stream_conv2d_2_source_37_pat_count_2 == 0)) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_3 <= _source_stream_conv2d_2_source_37_pat_cur_offset_3 + _source_stream_conv2d_2_source_37_pat_stride_buf_3;
        _source_stream_conv2d_2_source_37_pat_count_3 <= _source_stream_conv2d_2_source_37_pat_count_3 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_2_source_37_pat_count_0 == 0) && (_source_stream_conv2d_2_source_37_pat_count_1 == 0) && (_source_stream_conv2d_2_source_37_pat_count_2 == 0)) && (_source_stream_conv2d_2_source_37_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
        _source_stream_conv2d_2_source_37_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_2_source_37_pat_count_3 <= _source_stream_conv2d_2_source_37_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 1) && _stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_37_source_ram_renable <= 0;
        _stream_conv2d_2_source_37_idle <= 1;
      end 
      if((_stream_conv2d_2_source_37_source_pat_fsm_17 == 2) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_source_37_source_ram_renable <= 0;
        _stream_conv2d_2_source_37_idle <= 1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_251 <= _set_flag_250;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_252 <= _tmp_251;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_253 <= _tmp_252;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_254 <= _tmp_253;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_255 <= _tmp_254;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_256 <= _tmp_255;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_257 <= _tmp_256;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_258 <= _tmp_257;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_259 <= _tmp_258;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_260 <= _tmp_259;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_261 <= _tmp_260;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_262 <= _tmp_261;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_263 <= _tmp_262;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_264 <= _tmp_263;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_265 <= _tmp_264;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_266 <= _tmp_265;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_267 <= _tmp_266;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_268 <= _tmp_267;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_269 <= _tmp_268;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_270 <= _tmp_269;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_271 <= _tmp_270;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_272 <= _tmp_271;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_273 <= _tmp_272;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_274 <= _tmp_273;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_275 <= _tmp_274;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_276 <= _tmp_275;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_277 <= _tmp_276;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_278 <= _tmp_277;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_279 <= _tmp_278;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_280 <= _tmp_279;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_281 <= _tmp_280;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_284 <= _tmp_283;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_285 <= _tmp_284;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_286 <= _tmp_285;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_287 <= _tmp_286;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_288 <= _tmp_287;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_289 <= _tmp_288;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_290 <= _tmp_289;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_291 <= _tmp_290;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_292 <= _tmp_291;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_293 <= _tmp_292;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_294 <= _tmp_293;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_295 <= _tmp_294;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_296 <= _tmp_295;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_297 <= _tmp_296;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_298 <= _tmp_297;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_299 <= _tmp_298;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_300 <= _tmp_299;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_301 <= _tmp_300;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_302 <= _tmp_301;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_303 <= _tmp_302;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_304 <= _tmp_303;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_305 <= _tmp_304;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_306 <= _tmp_305;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_307 <= _tmp_306;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_308 <= _tmp_307;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_309 <= _tmp_308;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_310 <= _tmp_309;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_311 <= _tmp_310;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_312 <= _tmp_311;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_313 <= _tmp_312;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_314 <= _tmp_313;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_315 <= conv2d_2_next_stream_num_ops;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_316 <= _tmp_315;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_317 <= _tmp_316;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_318 <= _tmp_317;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_319 <= _tmp_318;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_320 <= _tmp_319;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_321 <= _tmp_320;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_322 <= _tmp_321;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_323 <= _tmp_322;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_324 <= _tmp_323;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_325 <= _tmp_324;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_326 <= _tmp_325;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_327 <= _tmp_326;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_328 <= _tmp_327;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_329 <= _tmp_328;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_330 <= _tmp_329;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_331 <= _tmp_330;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_332 <= _tmp_331;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_333 <= _tmp_332;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_334 <= _tmp_333;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_335 <= _tmp_334;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_336 <= _tmp_335;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_337 <= _tmp_336;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_338 <= _tmp_337;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_339 <= _tmp_338;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_340 <= _tmp_339;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_341 <= _tmp_340;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_342 <= _tmp_341;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_343 <= _tmp_342;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_344 <= _tmp_343;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_345 <= _tmp_344;
      end 
      if(_tmp_281) begin
        _stream_conv2d_2_sink_50_sink_mode <= 5'b1;
        _stream_conv2d_2_sink_50_sink_offset <= _tmp_314;
        _stream_conv2d_2_sink_50_sink_size <= _tmp_345;
        _stream_conv2d_2_sink_50_sink_stride <= 1;
      end 
      if(_tmp_281) begin
        _stream_conv2d_2_sink_50_sink_sel <= 19;
      end 
      if(_stream_conv2d_2_sink_start && _stream_conv2d_2_sink_50_sink_mode & 5'b1 && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_sink_50_sink_offset_buf <= _stream_conv2d_2_sink_50_sink_offset;
        _stream_conv2d_2_sink_50_sink_size_buf <= _stream_conv2d_2_sink_50_sink_size;
        _stream_conv2d_2_sink_50_sink_stride_buf <= _stream_conv2d_2_sink_50_sink_stride;
      end 
      if((_stream_conv2d_2_sink_50_sink_fsm_18 == 1) && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_sink_50_sink_waddr <= _stream_conv2d_2_sink_50_sink_offset_buf - _stream_conv2d_2_sink_50_sink_stride_buf;
        _stream_conv2d_2_sink_50_sink_count <= _stream_conv2d_2_sink_50_sink_size_buf;
      end 
      if((_stream_conv2d_2_sink_50_sink_fsm_18 == 2) && stream_conv2d_2_sink_51_data && _stream_conv2d_2_stream_oready) begin
        _stream_conv2d_2_sink_50_sink_waddr <= _stream_conv2d_2_sink_50_sink_waddr + _stream_conv2d_2_sink_50_sink_stride_buf;
        _stream_conv2d_2_sink_50_sink_wdata <= stream_conv2d_2_sink_50_data;
        _stream_conv2d_2_sink_50_sink_wenable <= 1;
        _stream_conv2d_2_sink_50_sink_count <= _stream_conv2d_2_sink_50_sink_count - 1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_735 <= _stream_conv2d_2_source_start;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_736 <= _tmp_735;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_737 <= _tmp_736;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_738 <= _stream_conv2d_2_source_start;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_739 <= _tmp_738;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_740 <= _tmp_739;
      end 
      if(_stream_conv2d_2_stream_oready && _tmp_740) begin
        __variable_wdata_264 <= 1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_741 <= _stream_conv2d_2_source_start;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_742 <= _tmp_741;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_743 <= _tmp_742;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_744 <= _tmp_743;
      end 
      if(_stream_conv2d_2_stream_oready && _tmp_744) begin
        __variable_wdata_264 <= 0;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_747 <= _tmp_746;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_750 <= _tmp_749;
      end 
      if(_stream_conv2d_2_stream_oready && _tmp_750) begin
        __variable_wdata_264 <= 1;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_751 <= _stream_conv2d_2_source_start;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_752 <= _tmp_751;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_753 <= _tmp_752;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_754 <= _tmp_753;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_755 <= _tmp_754;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_756 <= _tmp_755;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_757 <= _tmp_756;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_758 <= _tmp_757;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_759 <= _tmp_758;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_760 <= _tmp_759;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_761 <= _tmp_760;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_762 <= _tmp_761;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_763 <= _tmp_762;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_764 <= _tmp_763;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_765 <= _tmp_764;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_766 <= _tmp_765;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_767 <= _tmp_766;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_768 <= _tmp_767;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_769 <= _tmp_768;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_770 <= _tmp_769;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_771 <= _tmp_770;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_772 <= _tmp_771;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_773 <= _tmp_772;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_774 <= _tmp_773;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_775 <= _tmp_774;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_776 <= _tmp_775;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_777 <= _tmp_776;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_778 <= _tmp_777;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_779 <= _tmp_778;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_780 <= _tmp_779;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_781 <= _tmp_780;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_782 <= _stream_conv2d_2_source_stop;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_783 <= _tmp_782;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_784 <= _tmp_783;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_785 <= _tmp_784;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_786 <= _tmp_785;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_787 <= _tmp_786;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_788 <= _tmp_787;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_789 <= _tmp_788;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_790 <= _tmp_789;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_791 <= _tmp_790;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_792 <= _tmp_791;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_793 <= _tmp_792;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_794 <= _tmp_793;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_795 <= _tmp_794;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_796 <= _tmp_795;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_797 <= _tmp_796;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_798 <= _tmp_797;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_799 <= _tmp_798;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_800 <= _tmp_799;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_801 <= _tmp_800;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_802 <= _tmp_801;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_803 <= _tmp_802;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_804 <= _tmp_803;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_805 <= _tmp_804;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_806 <= _tmp_805;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_807 <= _tmp_806;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_808 <= _tmp_807;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_809 <= _tmp_808;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_810 <= _tmp_809;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_811 <= _tmp_810;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_812 <= _tmp_811;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_813 <= _stream_conv2d_2_source_busy;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_814 <= _tmp_813;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_815 <= _tmp_814;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_816 <= _tmp_815;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_817 <= _tmp_816;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_818 <= _tmp_817;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_819 <= _tmp_818;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_820 <= _tmp_819;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_821 <= _tmp_820;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_822 <= _tmp_821;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_823 <= _tmp_822;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_824 <= _tmp_823;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_825 <= _tmp_824;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_826 <= _tmp_825;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_827 <= _tmp_826;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_828 <= _tmp_827;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_829 <= _tmp_828;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_830 <= _tmp_829;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_831 <= _tmp_830;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_832 <= _tmp_831;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_833 <= _tmp_832;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_834 <= _tmp_833;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_835 <= _tmp_834;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_836 <= _tmp_835;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_837 <= _tmp_836;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_838 <= _tmp_837;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_839 <= _tmp_838;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_840 <= _tmp_839;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_841 <= _tmp_840;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_842 <= _tmp_841;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_843 <= _tmp_842;
      end 
      if(_stream_conv2d_2_stream_oready) begin
        _tmp_844 <= _stream_conv2d_2_sink_busy;
      end 
      if(!_stream_conv2d_2_sink_busy && _tmp_844) begin
        _stream_conv2d_2_busy_reg <= 0;
      end 
      if(_stream_conv2d_2_source_busy) begin
        _stream_conv2d_2_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_conv2d_2_fsm_1 = 1;
  localparam _stream_conv2d_2_fsm_2 = 2;
  localparam _stream_conv2d_2_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_fsm <= _stream_conv2d_2_fsm_init;
      _stream_conv2d_2_source_start <= 0;
      _stream_conv2d_2_source_busy <= 0;
      _stream_conv2d_2_stream_ivalid <= 0;
    end else begin
      if(_stream_conv2d_2_stream_oready && _tmp_737) begin
        _stream_conv2d_2_stream_ivalid <= 1;
      end 
      if(_stream_conv2d_2_stream_oready && _tmp_747) begin
        _stream_conv2d_2_stream_ivalid <= 0;
      end 
      case(_stream_conv2d_2_fsm)
        _stream_conv2d_2_fsm_init: begin
          if(_stream_conv2d_2_run_flag) begin
            _stream_conv2d_2_source_start <= 1;
          end 
          if(_stream_conv2d_2_run_flag) begin
            _stream_conv2d_2_fsm <= _stream_conv2d_2_fsm_1;
          end 
        end
        _stream_conv2d_2_fsm_1: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_start <= 0;
            _stream_conv2d_2_source_busy <= 1;
          end 
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_fsm <= _stream_conv2d_2_fsm_2;
          end 
        end
        _stream_conv2d_2_fsm_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_fsm <= _stream_conv2d_2_fsm_3;
          end 
        end
        _stream_conv2d_2_fsm_3: begin
          if(_stream_conv2d_2_stream_oready && (_stream_conv2d_2_source_11_idle && _stream_conv2d_2_source_13_idle && _stream_conv2d_2_source_15_idle && _stream_conv2d_2_source_20_idle && _stream_conv2d_2_source_21_idle && _stream_conv2d_2_source_22_idle && _stream_conv2d_2_source_23_idle && _stream_conv2d_2_source_24_idle && _stream_conv2d_2_source_25_idle && _stream_conv2d_2_source_26_idle && _stream_conv2d_2_source_27_idle && _stream_conv2d_2_source_28_idle && _stream_conv2d_2_source_29_idle && _stream_conv2d_2_source_30_idle && _stream_conv2d_2_source_31_idle && _stream_conv2d_2_source_32_idle && _stream_conv2d_2_source_33_idle && _stream_conv2d_2_source_34_idle && _stream_conv2d_2_source_35_idle && _stream_conv2d_2_source_36_idle && _stream_conv2d_2_source_37_idle && _stream_conv2d_2_source_7_idle && _stream_conv2d_2_source_9_idle && (_stream_conv2d_2_fsm == 3))) begin
            _stream_conv2d_2_source_busy <= 0;
          end 
          if(_stream_conv2d_2_stream_oready && (_stream_conv2d_2_source_11_idle && _stream_conv2d_2_source_13_idle && _stream_conv2d_2_source_15_idle && _stream_conv2d_2_source_20_idle && _stream_conv2d_2_source_21_idle && _stream_conv2d_2_source_22_idle && _stream_conv2d_2_source_23_idle && _stream_conv2d_2_source_24_idle && _stream_conv2d_2_source_25_idle && _stream_conv2d_2_source_26_idle && _stream_conv2d_2_source_27_idle && _stream_conv2d_2_source_28_idle && _stream_conv2d_2_source_29_idle && _stream_conv2d_2_source_30_idle && _stream_conv2d_2_source_31_idle && _stream_conv2d_2_source_32_idle && _stream_conv2d_2_source_33_idle && _stream_conv2d_2_source_34_idle && _stream_conv2d_2_source_35_idle && _stream_conv2d_2_source_36_idle && _stream_conv2d_2_source_37_idle && _stream_conv2d_2_source_7_idle && _stream_conv2d_2_source_9_idle && (_stream_conv2d_2_fsm == 3)) && _stream_conv2d_2_run_flag) begin
            _stream_conv2d_2_source_start <= 1;
          end 
          if(_stream_conv2d_2_stream_oready && (_stream_conv2d_2_source_11_idle && _stream_conv2d_2_source_13_idle && _stream_conv2d_2_source_15_idle && _stream_conv2d_2_source_20_idle && _stream_conv2d_2_source_21_idle && _stream_conv2d_2_source_22_idle && _stream_conv2d_2_source_23_idle && _stream_conv2d_2_source_24_idle && _stream_conv2d_2_source_25_idle && _stream_conv2d_2_source_26_idle && _stream_conv2d_2_source_27_idle && _stream_conv2d_2_source_28_idle && _stream_conv2d_2_source_29_idle && _stream_conv2d_2_source_30_idle && _stream_conv2d_2_source_31_idle && _stream_conv2d_2_source_32_idle && _stream_conv2d_2_source_33_idle && _stream_conv2d_2_source_34_idle && _stream_conv2d_2_source_35_idle && _stream_conv2d_2_source_36_idle && _stream_conv2d_2_source_37_idle && _stream_conv2d_2_source_7_idle && _stream_conv2d_2_source_9_idle && (_stream_conv2d_2_fsm == 3))) begin
            _stream_conv2d_2_fsm <= _stream_conv2d_2_fsm_init;
          end 
          if(_stream_conv2d_2_stream_oready && (_stream_conv2d_2_source_11_idle && _stream_conv2d_2_source_13_idle && _stream_conv2d_2_source_15_idle && _stream_conv2d_2_source_20_idle && _stream_conv2d_2_source_21_idle && _stream_conv2d_2_source_22_idle && _stream_conv2d_2_source_23_idle && _stream_conv2d_2_source_24_idle && _stream_conv2d_2_source_25_idle && _stream_conv2d_2_source_26_idle && _stream_conv2d_2_source_27_idle && _stream_conv2d_2_source_28_idle && _stream_conv2d_2_source_29_idle && _stream_conv2d_2_source_30_idle && _stream_conv2d_2_source_31_idle && _stream_conv2d_2_source_32_idle && _stream_conv2d_2_source_33_idle && _stream_conv2d_2_source_34_idle && _stream_conv2d_2_source_35_idle && _stream_conv2d_2_source_36_idle && _stream_conv2d_2_source_37_idle && _stream_conv2d_2_source_7_idle && _stream_conv2d_2_source_9_idle && (_stream_conv2d_2_fsm == 3)) && _stream_conv2d_2_run_flag) begin
            _stream_conv2d_2_fsm <= _stream_conv2d_2_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_celu_3_source_1_source_ram_renable <= 0;
      _stream_celu_3_source_1_source_fifo_deq <= 0;
      _stream_celu_3_source_1_idle <= 1;
      _stream_celu_3_sink_2_sink_wenable <= 0;
      _stream_celu_3_sink_2_sink_fifo_enq <= 0;
      __stream_celu_3_stream_ivalid_1 <= 0;
      __stream_celu_3_stream_ivalid_2 <= 0;
      __stream_celu_3_stream_ivalid_3 <= 0;
      __stream_celu_3_stream_ivalid_4 <= 0;
      __stream_celu_3_stream_ivalid_5 <= 0;
      __stream_celu_3_stream_ivalid_6 <= 0;
      __stream_celu_3_stream_ivalid_7 <= 0;
      __stream_celu_3_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_849 <= 0;
      _greatereq_data_862 <= 0;
      __delay_data_999_reinterpretcast_850 <= 0;
      __delay_data_1009_reinterpretcast_846 <= 0;
      __delay_data_1000__delay_999_reinterpretcast_850 <= 0;
      __delay_data_1003_greatereq_862 <= 0;
      __delay_data_1010__delay_1009_reinterpretcast_846 <= 0;
      __delay_data_1001__delay_1000__delay_999_reinterpretcast_850 <= 0;
      __delay_data_1004__delay_1003_greatereq_862 <= 0;
      __delay_data_1011__delay_1010__delay_1009_reinterpretcast_846 <= 0;
      _abs_data_852 <= 0;
      __delay_data_1002__delay_1001__delay_1000___reinterpretcast_850 <= 0;
      __delay_data_1005__delay_1004__delay_1003_greatereq_862 <= 0;
      __delay_data_1012__delay_1011__delay_1010___reinterpretcast_846 <= 0;
      _sra_data_853 <= 0;
      __delay_data_1006__delay_1005__delay_1004___greatereq_862 <= 0;
      __delay_data_1013__delay_1012__delay_1011___reinterpretcast_846 <= 0;
      _greaterthan_data_858 <= 0;
      __delay_data_1007__delay_1006__delay_1005___greatereq_862 <= 0;
      __delay_data_1014__delay_1013__delay_1012___reinterpretcast_846 <= 0;
      _cond_data_860 <= 0;
      __delay_data_1008__delay_1007__delay_1006___greatereq_862 <= 0;
      __delay_data_1015__delay_1014__delay_1013___reinterpretcast_846 <= 0;
      _cond_data_864 <= 0;
      _stream_celu_3_parameter_0_next_parameter_data <= 0;
      __variable_wdata_844 <= 0;
      _stream_celu_3_source_1_source_mode <= 5'b0;
      _stream_celu_3_source_1_source_offset <= 0;
      _stream_celu_3_source_1_source_size <= 0;
      _stream_celu_3_source_1_source_stride <= 0;
      _stream_celu_3_source_1_source_sel <= 0;
      _stream_celu_3_source_1_source_offset_buf <= 0;
      _stream_celu_3_source_1_source_size_buf <= 0;
      _stream_celu_3_source_1_source_stride_buf <= 0;
      __variable_wdata_845 <= 0;
      _stream_celu_3_source_1_source_ram_raddr <= 0;
      _stream_celu_3_source_1_source_count <= 0;
      _tmp_896 <= 0;
      _tmp_897 <= 0;
      _tmp_898 <= 0;
      _tmp_899 <= 0;
      _tmp_900 <= 0;
      _tmp_901 <= 0;
      _tmp_902 <= 0;
      _tmp_903 <= 0;
      _tmp_904 <= 0;
      _tmp_905 <= 0;
      _tmp_906 <= 0;
      _tmp_907 <= 0;
      _tmp_908 <= 0;
      _tmp_909 <= 0;
      _tmp_910 <= 0;
      _tmp_911 <= 0;
      _tmp_912 <= 0;
      _tmp_913 <= 0;
      _tmp_914 <= 0;
      _tmp_915 <= 0;
      _tmp_916 <= 0;
      _tmp_917 <= 0;
      _tmp_918 <= 0;
      _tmp_919 <= 0;
      _tmp_920 <= 0;
      _tmp_921 <= 0;
      _tmp_922 <= 0;
      _tmp_923 <= 0;
      _tmp_924 <= 0;
      _tmp_925 <= 0;
      _stream_celu_3_sink_2_sink_mode <= 5'b0;
      _stream_celu_3_sink_2_sink_offset <= 0;
      _stream_celu_3_sink_2_sink_size <= 0;
      _stream_celu_3_sink_2_sink_stride <= 0;
      _stream_celu_3_sink_2_sink_sel <= 0;
      _stream_celu_3_sink_2_sink_offset_buf <= 0;
      _stream_celu_3_sink_2_sink_size_buf <= 0;
      _stream_celu_3_sink_2_sink_stride_buf <= 0;
      _stream_celu_3_sink_2_sink_waddr <= 0;
      _stream_celu_3_sink_2_sink_count <= 0;
      _stream_celu_3_sink_2_sink_wdata <= 0;
      _tmp_927 <= 0;
      _tmp_928 <= 0;
      _tmp_929 <= 0;
      _tmp_932 <= 0;
      _tmp_933 <= 0;
      _tmp_934 <= 0;
      _tmp_935 <= 0;
      _tmp_936 <= 0;
      _tmp_937 <= 0;
      _tmp_938 <= 0;
      _tmp_939 <= 0;
      _tmp_940 <= 0;
      _tmp_941 <= 0;
      _tmp_942 <= 0;
      _tmp_943 <= 0;
      _tmp_944 <= 0;
      _tmp_945 <= 0;
      _tmp_946 <= 0;
      _tmp_947 <= 0;
      _tmp_948 <= 0;
      _tmp_949 <= 0;
      _tmp_950 <= 0;
      _tmp_951 <= 0;
      _tmp_952 <= 0;
      _tmp_953 <= 0;
      _tmp_954 <= 0;
      _tmp_955 <= 0;
      _tmp_956 <= 0;
      _tmp_957 <= 0;
      _tmp_958 <= 0;
      _tmp_959 <= 0;
      _tmp_960 <= 0;
      _tmp_961 <= 0;
      _tmp_962 <= 0;
      _tmp_963 <= 0;
      _stream_celu_3_busy_reg <= 0;
    end else begin
      if(_stream_celu_3_stream_oready) begin
        _stream_celu_3_source_1_source_ram_renable <= 0;
        _stream_celu_3_source_1_source_fifo_deq <= 0;
      end 
      _stream_celu_3_source_1_idle <= _stream_celu_3_source_1_idle;
      if(_stream_celu_3_stream_oready) begin
        _stream_celu_3_sink_2_sink_wenable <= 0;
        _stream_celu_3_sink_2_sink_fifo_enq <= 0;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_1 <= _stream_celu_3_stream_ivalid;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_2 <= __stream_celu_3_stream_ivalid_1;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_3 <= __stream_celu_3_stream_ivalid_2;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_4 <= __stream_celu_3_stream_ivalid_3;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_5 <= __stream_celu_3_stream_ivalid_4;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_6 <= __stream_celu_3_stream_ivalid_5;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_7 <= __stream_celu_3_stream_ivalid_6;
      end 
      if(_stream_celu_3_stream_oready) begin
        __stream_celu_3_stream_ivalid_8 <= __stream_celu_3_stream_ivalid_7;
      end 
      if(_stream_celu_3_stream_oready) begin
        _times_mul_odata_reg_849 <= _times_mul_odata_849;
      end 
      if(_stream_celu_3_stream_oready) begin
        _greatereq_data_862 <= _reinterpretcast_data_846 >= 1'sd0;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_999_reinterpretcast_850 <= _reinterpretcast_data_850;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1009_reinterpretcast_846 <= _reinterpretcast_data_846;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1000__delay_999_reinterpretcast_850 <= __delay_data_999_reinterpretcast_850;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1003_greatereq_862 <= _greatereq_data_862;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1010__delay_1009_reinterpretcast_846 <= __delay_data_1009_reinterpretcast_846;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1001__delay_1000__delay_999_reinterpretcast_850 <= __delay_data_1000__delay_999_reinterpretcast_850;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1004__delay_1003_greatereq_862 <= __delay_data_1003_greatereq_862;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1011__delay_1010__delay_1009_reinterpretcast_846 <= __delay_data_1010__delay_1009_reinterpretcast_846;
      end 
      if(_stream_celu_3_stream_oready) begin
        _abs_data_852 <= (_times_data_849 < 'sd0)? ~_times_data_849 + 1 : _times_data_849;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1002__delay_1001__delay_1000___reinterpretcast_850 <= __delay_data_1001__delay_1000__delay_999_reinterpretcast_850;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1005__delay_1004__delay_1003_greatereq_862 <= __delay_data_1004__delay_1003_greatereq_862;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1012__delay_1011__delay_1010___reinterpretcast_846 <= __delay_data_1011__delay_1010__delay_1009_reinterpretcast_846;
      end 
      if(_stream_celu_3_stream_oready) begin
        _sra_data_853 <= _abs_data_852 >>> __delay_data_1002__delay_1001__delay_1000___reinterpretcast_850;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1006__delay_1005__delay_1004___greatereq_862 <= __delay_data_1005__delay_1004__delay_1003_greatereq_862;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1013__delay_1012__delay_1011___reinterpretcast_846 <= __delay_data_1012__delay_1011__delay_1010___reinterpretcast_846;
      end 
      if(_stream_celu_3_stream_oready) begin
        _greaterthan_data_858 <= _sra_data_853 > 9'sd255;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1007__delay_1006__delay_1005___greatereq_862 <= __delay_data_1006__delay_1005__delay_1004___greatereq_862;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1014__delay_1013__delay_1012___reinterpretcast_846 <= __delay_data_1013__delay_1012__delay_1011___reinterpretcast_846;
      end 
      if(_stream_celu_3_stream_oready) begin
        _cond_data_860 <= (_greaterthan_data_858)? -33'sd2147483648 : _lut_data_857;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1008__delay_1007__delay_1006___greatereq_862 <= __delay_data_1007__delay_1006__delay_1005___greatereq_862;
      end 
      if(_stream_celu_3_stream_oready) begin
        __delay_data_1015__delay_1014__delay_1013___reinterpretcast_846 <= __delay_data_1014__delay_1013__delay_1012___reinterpretcast_846;
      end 
      if(_stream_celu_3_stream_oready) begin
        _cond_data_864 <= (__delay_data_1008__delay_1007__delay_1006___greatereq_862)? __delay_data_1015__delay_1014__delay_1013___reinterpretcast_846 : _cond_data_860;
      end 
      if(_set_flag_891) begin
        _stream_celu_3_parameter_0_next_parameter_data <= (cparam_celu_3_arg_stride_zeros_0)? 1 : 0;
      end 
      if(_stream_celu_3_source_start) begin
        __variable_wdata_844 <= _stream_celu_3_parameter_0_next_parameter_data;
      end 
      if(_set_flag_892) begin
        _stream_celu_3_source_1_source_mode <= 5'b1;
        _stream_celu_3_source_1_source_offset <= celu_3_arg_page_comp_offset_0;
        _stream_celu_3_source_1_source_size <= cparam_celu_3_dma_size;
        _stream_celu_3_source_1_source_stride <= (cparam_celu_3_arg_stride_zeros_0)? 0 : 1;
      end 
      if(_set_flag_892) begin
        _stream_celu_3_source_1_source_sel <= 1;
      end 
      if(_stream_celu_3_source_start && _stream_celu_3_source_1_source_mode & 5'b1 && _stream_celu_3_stream_oready) begin
        _stream_celu_3_source_1_source_offset_buf <= _stream_celu_3_source_1_source_offset;
        _stream_celu_3_source_1_source_size_buf <= _stream_celu_3_source_1_source_size;
        _stream_celu_3_source_1_source_stride_buf <= _stream_celu_3_source_1_source_stride;
      end 
      if(_stream_celu_3_stream_oready && _stream_celu_3_source_busy && _stream_celu_3_is_root) begin
        __variable_wdata_845 <= _stream_celu_3_source_1_source_ram_rdata;
      end 
      if((_stream_celu_3_source_1_source_fsm_0 == 1) && _stream_celu_3_stream_oready) begin
        _stream_celu_3_source_1_idle <= 0;
        _stream_celu_3_source_1_source_ram_raddr <= _stream_celu_3_source_1_source_offset_buf;
        _stream_celu_3_source_1_source_ram_renable <= 1;
        _stream_celu_3_source_1_source_count <= _stream_celu_3_source_1_source_size_buf;
      end 
      if((_stream_celu_3_source_1_source_fsm_0 == 2) && _stream_celu_3_stream_oready) begin
        _stream_celu_3_source_1_source_ram_raddr <= _stream_celu_3_source_1_source_ram_raddr + _stream_celu_3_source_1_source_stride_buf;
        _stream_celu_3_source_1_source_ram_renable <= 1;
        _stream_celu_3_source_1_source_count <= _stream_celu_3_source_1_source_count - 1;
      end 
      if((_stream_celu_3_source_1_source_fsm_0 == 2) && (_stream_celu_3_source_1_source_count == 1) && _stream_celu_3_stream_oready) begin
        _stream_celu_3_source_1_source_ram_renable <= 0;
        _stream_celu_3_source_1_idle <= 1;
      end 
      if((_stream_celu_3_source_1_source_fsm_0 == 2) && _stream_celu_3_source_stop && _stream_celu_3_stream_oready) begin
        _stream_celu_3_source_1_source_ram_renable <= 0;
        _stream_celu_3_source_1_idle <= 1;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_896 <= _set_flag_895;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_897 <= _tmp_896;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_898 <= _tmp_897;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_899 <= _tmp_898;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_900 <= _tmp_899;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_901 <= _tmp_900;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_902 <= _tmp_901;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_903 <= _tmp_902;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_904 <= _tmp_903;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_905 <= _tmp_904;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_906 <= celu_3_out_page_comp_offset;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_907 <= _tmp_906;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_908 <= _tmp_907;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_909 <= _tmp_908;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_910 <= _tmp_909;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_911 <= _tmp_910;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_912 <= _tmp_911;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_913 <= _tmp_912;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_914 <= _tmp_913;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_915 <= _tmp_914;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_916 <= cparam_celu_3_dma_size;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_917 <= _tmp_916;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_918 <= _tmp_917;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_919 <= _tmp_918;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_920 <= _tmp_919;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_921 <= _tmp_920;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_922 <= _tmp_921;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_923 <= _tmp_922;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_924 <= _tmp_923;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_925 <= _tmp_924;
      end 
      if(_tmp_905) begin
        _stream_celu_3_sink_2_sink_mode <= 5'b1;
        _stream_celu_3_sink_2_sink_offset <= _tmp_915;
        _stream_celu_3_sink_2_sink_size <= _tmp_925;
        _stream_celu_3_sink_2_sink_stride <= 1;
      end 
      if(_tmp_905) begin
        _stream_celu_3_sink_2_sink_sel <= 2;
      end 
      if(_stream_celu_3_sink_start && _stream_celu_3_sink_2_sink_mode & 5'b1 && _stream_celu_3_stream_oready) begin
        _stream_celu_3_sink_2_sink_offset_buf <= _stream_celu_3_sink_2_sink_offset;
        _stream_celu_3_sink_2_sink_size_buf <= _stream_celu_3_sink_2_sink_size;
        _stream_celu_3_sink_2_sink_stride_buf <= _stream_celu_3_sink_2_sink_stride;
      end 
      if((_stream_celu_3_sink_2_sink_fsm_1 == 1) && _stream_celu_3_stream_oready) begin
        _stream_celu_3_sink_2_sink_waddr <= _stream_celu_3_sink_2_sink_offset_buf - _stream_celu_3_sink_2_sink_stride_buf;
        _stream_celu_3_sink_2_sink_count <= _stream_celu_3_sink_2_sink_size_buf;
      end 
      if((_stream_celu_3_sink_2_sink_fsm_1 == 2) && _stream_celu_3_stream_oready) begin
        _stream_celu_3_sink_2_sink_waddr <= _stream_celu_3_sink_2_sink_waddr + _stream_celu_3_sink_2_sink_stride_buf;
        _stream_celu_3_sink_2_sink_wdata <= stream_celu_3_sink_2_data;
        _stream_celu_3_sink_2_sink_wenable <= 1;
        _stream_celu_3_sink_2_sink_count <= _stream_celu_3_sink_2_sink_count - 1;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_927 <= _stream_celu_3_source_start;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_928 <= _tmp_927;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_929 <= _tmp_928;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_932 <= _tmp_931;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_933 <= _stream_celu_3_source_start;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_934 <= _tmp_933;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_935 <= _tmp_934;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_936 <= _tmp_935;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_937 <= _tmp_936;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_938 <= _tmp_937;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_939 <= _tmp_938;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_940 <= _tmp_939;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_941 <= _tmp_940;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_942 <= _tmp_941;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_943 <= _stream_celu_3_source_stop;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_944 <= _tmp_943;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_945 <= _tmp_944;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_946 <= _tmp_945;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_947 <= _tmp_946;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_948 <= _tmp_947;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_949 <= _tmp_948;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_950 <= _tmp_949;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_951 <= _tmp_950;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_952 <= _tmp_951;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_953 <= _stream_celu_3_source_busy;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_954 <= _tmp_953;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_955 <= _tmp_954;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_956 <= _tmp_955;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_957 <= _tmp_956;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_958 <= _tmp_957;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_959 <= _tmp_958;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_960 <= _tmp_959;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_961 <= _tmp_960;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_962 <= _tmp_961;
      end 
      if(_stream_celu_3_stream_oready) begin
        _tmp_963 <= _stream_celu_3_sink_busy;
      end 
      if(!_stream_celu_3_sink_busy && _tmp_963) begin
        _stream_celu_3_busy_reg <= 0;
      end 
      if(_stream_celu_3_source_busy) begin
        _stream_celu_3_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_celu_3_fsm_1 = 1;
  localparam _stream_celu_3_fsm_2 = 2;
  localparam _stream_celu_3_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_celu_3_fsm <= _stream_celu_3_fsm_init;
      _stream_celu_3_source_start <= 0;
      _stream_celu_3_source_busy <= 0;
      _stream_celu_3_stream_ivalid <= 0;
    end else begin
      if(_stream_celu_3_stream_oready && _tmp_929) begin
        _stream_celu_3_stream_ivalid <= 1;
      end 
      if(_stream_celu_3_stream_oready && _tmp_932) begin
        _stream_celu_3_stream_ivalid <= 0;
      end 
      case(_stream_celu_3_fsm)
        _stream_celu_3_fsm_init: begin
          if(_stream_celu_3_run_flag) begin
            _stream_celu_3_source_start <= 1;
          end 
          if(_stream_celu_3_run_flag) begin
            _stream_celu_3_fsm <= _stream_celu_3_fsm_1;
          end 
        end
        _stream_celu_3_fsm_1: begin
          if(_stream_celu_3_source_start && _stream_celu_3_stream_oready) begin
            _stream_celu_3_source_start <= 0;
            _stream_celu_3_source_busy <= 1;
          end 
          if(_stream_celu_3_source_start && _stream_celu_3_stream_oready) begin
            _stream_celu_3_fsm <= _stream_celu_3_fsm_2;
          end 
        end
        _stream_celu_3_fsm_2: begin
          if(_stream_celu_3_stream_oready) begin
            _stream_celu_3_fsm <= _stream_celu_3_fsm_3;
          end 
        end
        _stream_celu_3_fsm_3: begin
          if(_stream_celu_3_stream_oready && (_stream_celu_3_source_1_idle && (_stream_celu_3_fsm == 3))) begin
            _stream_celu_3_source_busy <= 0;
          end 
          if(_stream_celu_3_stream_oready && (_stream_celu_3_source_1_idle && (_stream_celu_3_fsm == 3)) && _stream_celu_3_run_flag) begin
            _stream_celu_3_source_start <= 1;
          end 
          if(_stream_celu_3_stream_oready && (_stream_celu_3_source_1_idle && (_stream_celu_3_fsm == 3))) begin
            _stream_celu_3_fsm <= _stream_celu_3_fsm_init;
          end 
          if(_stream_celu_3_stream_oready && (_stream_celu_3_source_1_idle && (_stream_celu_3_fsm == 3)) && _stream_celu_3_run_flag) begin
            _stream_celu_3_fsm <= _stream_celu_3_fsm_1;
          end 
        end
      endcase
    end
  end

  localparam main_fsm_1 = 1;
  localparam main_fsm_2 = 2;
  localparam main_fsm_3 = 3;
  localparam main_fsm_4 = 4;
  localparam main_fsm_5 = 5;
  localparam main_fsm_6 = 6;
  localparam main_fsm_7 = 7;
  localparam main_fsm_8 = 8;
  localparam main_fsm_9 = 9;
  localparam main_fsm_10 = 10;
  localparam main_fsm_11 = 11;
  localparam main_fsm_12 = 12;
  localparam main_fsm_13 = 13;
  localparam main_fsm_14 = 14;
  localparam main_fsm_15 = 15;
  localparam main_fsm_16 = 16;
  localparam main_fsm_17 = 17;
  localparam main_fsm_18 = 18;
  localparam main_fsm_19 = 19;
  localparam main_fsm_20 = 20;
  localparam main_fsm_21 = 21;
  localparam main_fsm_22 = 22;

  always @(posedge CLK) begin
    if(RST) begin
      main_fsm <= main_fsm_init;
      conv2d_2_objaddr <= 0;
      conv2d_2_arg_objaddr_0 <= 0;
      conv2d_2_arg_objaddr_1 <= 0;
      celu_3_objaddr <= 0;
      celu_3_arg_objaddr_0 <= 0;
    end else begin
      case(main_fsm)
        main_fsm_init: begin
          if(_saxi_register_4 != 0) begin
            main_fsm <= main_fsm_1;
          end 
        end
        main_fsm_1: begin
          main_fsm <= main_fsm_2;
        end
        main_fsm_2: begin
          main_fsm <= main_fsm_3;
        end
        main_fsm_3: begin
          main_fsm <= main_fsm_4;
        end
        main_fsm_4: begin
          main_fsm <= main_fsm_5;
        end
        main_fsm_5: begin
          conv2d_2_objaddr <= _saxi_register_33;
          main_fsm <= main_fsm_6;
        end
        main_fsm_6: begin
          conv2d_2_arg_objaddr_0 <= _saxi_register_35;
          main_fsm <= main_fsm_7;
        end
        main_fsm_7: begin
          conv2d_2_arg_objaddr_1 <= _saxi_register_36;
          main_fsm <= main_fsm_8;
        end
        main_fsm_8: begin
          main_fsm <= main_fsm_9;
        end
        main_fsm_9: begin
          main_fsm <= main_fsm_10;
        end
        main_fsm_10: begin
          if(control_conv2d_2 == 30) begin
            main_fsm <= main_fsm_11;
          end 
        end
        main_fsm_11: begin
          main_fsm <= main_fsm_12;
        end
        main_fsm_12: begin
          celu_3_objaddr <= _saxi_register_34;
          main_fsm <= main_fsm_13;
        end
        main_fsm_13: begin
          celu_3_arg_objaddr_0 <= _saxi_register_33;
          main_fsm <= main_fsm_14;
        end
        main_fsm_14: begin
          main_fsm <= main_fsm_15;
        end
        main_fsm_15: begin
          main_fsm <= main_fsm_16;
        end
        main_fsm_16: begin
          if(control_celu_3 == 23) begin
            main_fsm <= main_fsm_17;
          end 
        end
        main_fsm_17: begin
          main_fsm <= main_fsm_18;
        end
        main_fsm_18: begin
          main_fsm <= main_fsm_19;
        end
        main_fsm_19: begin
          main_fsm <= main_fsm_20;
        end
        main_fsm_20: begin
          main_fsm <= main_fsm_21;
        end
        main_fsm_21: begin
          main_fsm <= main_fsm_22;
        end
        main_fsm_22: begin
          main_fsm <= main_fsm_init;
        end
      endcase
    end
  end

  localparam control_conv2d_2_1 = 1;
  localparam control_conv2d_2_2 = 2;
  localparam control_conv2d_2_3 = 3;
  localparam control_conv2d_2_4 = 4;
  localparam control_conv2d_2_5 = 5;
  localparam control_conv2d_2_6 = 6;
  localparam control_conv2d_2_7 = 7;
  localparam control_conv2d_2_8 = 8;
  localparam control_conv2d_2_9 = 9;
  localparam control_conv2d_2_10 = 10;
  localparam control_conv2d_2_11 = 11;
  localparam control_conv2d_2_12 = 12;
  localparam control_conv2d_2_13 = 13;
  localparam control_conv2d_2_14 = 14;
  localparam control_conv2d_2_15 = 15;
  localparam control_conv2d_2_16 = 16;
  localparam control_conv2d_2_17 = 17;
  localparam control_conv2d_2_18 = 18;
  localparam control_conv2d_2_19 = 19;
  localparam control_conv2d_2_20 = 20;
  localparam control_conv2d_2_21 = 21;
  localparam control_conv2d_2_22 = 22;
  localparam control_conv2d_2_23 = 23;
  localparam control_conv2d_2_24 = 24;
  localparam control_conv2d_2_25 = 25;
  localparam control_conv2d_2_26 = 26;
  localparam control_conv2d_2_27 = 27;
  localparam control_conv2d_2_28 = 28;
  localparam control_conv2d_2_29 = 29;
  localparam control_conv2d_2_30 = 30;

  always @(posedge CLK) begin
    if(RST) begin
      control_conv2d_2 <= control_conv2d_2_init;
      _control_conv2d_2_called <= 0;
      conv2d_2_filter_base_offset <= 0;
      conv2d_2_filter_page_comp_offset <= 0;
      conv2d_2_filter_page_dma_offset <= 0;
      conv2d_2_act_base_offset_row <= 0;
      conv2d_2_act_base_offset_bat <= 0;
      conv2d_2_dma_flag_0 <= 0;
      conv2d_2_dma_flag_1 <= 0;
      conv2d_2_dma_flag_2 <= 0;
      conv2d_2_act_page_comp_offset_0 <= 0;
      conv2d_2_act_page_comp_offset_1 <= 0;
      conv2d_2_act_page_comp_offset_2 <= 0;
      conv2d_2_act_page_dma_offset_0 <= 0;
      conv2d_2_act_page_dma_offset_1 <= 0;
      conv2d_2_act_page_dma_offset_2 <= 0;
      conv2d_2_out_base_offset_val <= 0;
      conv2d_2_out_base_offset_col <= 0;
      conv2d_2_out_base_offset_row <= 0;
      conv2d_2_out_base_offset_bat <= 0;
      conv2d_2_out_base_offset_och <= 0;
      conv2d_2_out_page <= 0;
      conv2d_2_out_page_comp_offset <= 0;
      conv2d_2_out_page_dma_offset <= 0;
      conv2d_2_out_laddr_offset <= 0;
      conv2d_2_sync_out_count <= 0;
      conv2d_2_write_count <= 0;
      conv2d_2_next_out_write_size <= 0;
      conv2d_2_row_count <= 0;
      conv2d_2_bat_count <= 0;
      conv2d_2_och_count <= 0;
      conv2d_2_row_select <= 0;
      conv2d_2_prev_row_count <= 0;
      conv2d_2_prev_bat_count <= 0;
      conv2d_2_prev_och_count <= 0;
      conv2d_2_prev_row_select <= 0;
      conv2d_2_out_col_count <= 0;
      conv2d_2_out_row_count <= 0;
      conv2d_2_out_ram_select <= 0;
      conv2d_2_skip_read_filter <= 0;
      conv2d_2_skip_read_act <= 0;
      conv2d_2_skip_comp <= 0;
      conv2d_2_skip_write_out <= 1;
    end else begin
      case(control_conv2d_2)
        control_conv2d_2_init: begin
          if(main_fsm == 8) begin
            _control_conv2d_2_called <= 1;
          end 
          if(main_fsm == 8) begin
            control_conv2d_2 <= control_conv2d_2_1;
          end 
        end
        control_conv2d_2_1: begin
          control_conv2d_2 <= control_conv2d_2_2;
        end
        control_conv2d_2_2: begin
          conv2d_2_filter_base_offset <= 0;
          conv2d_2_filter_page_comp_offset <= 0;
          conv2d_2_filter_page_dma_offset <= 0;
          conv2d_2_act_base_offset_row <= 0;
          conv2d_2_act_base_offset_bat <= 0;
          conv2d_2_dma_flag_0 <= 1;
          conv2d_2_dma_flag_1 <= 1;
          conv2d_2_dma_flag_2 <= 1;
          conv2d_2_act_page_comp_offset_0 <= 0;
          conv2d_2_act_page_comp_offset_1 <= 0;
          conv2d_2_act_page_comp_offset_2 <= 0;
          conv2d_2_act_page_dma_offset_0 <= 0;
          conv2d_2_act_page_dma_offset_1 <= 0;
          conv2d_2_act_page_dma_offset_2 <= 0;
          conv2d_2_out_base_offset_val <= 0;
          conv2d_2_out_base_offset_col <= 0;
          conv2d_2_out_base_offset_row <= 0;
          conv2d_2_out_base_offset_bat <= 0;
          conv2d_2_out_base_offset_och <= 0;
          conv2d_2_out_page <= 0;
          conv2d_2_out_page_comp_offset <= 0;
          conv2d_2_out_page_dma_offset <= 0;
          conv2d_2_out_laddr_offset <= 0;
          conv2d_2_sync_out_count <= 0;
          conv2d_2_write_count <= 0;
          conv2d_2_next_out_write_size <= (cparam_conv2d_2_max_och_count == 0)? cparam_conv2d_2_out_write_size_res : cparam_conv2d_2_out_write_size;
          conv2d_2_row_count <= 0;
          conv2d_2_bat_count <= 0;
          conv2d_2_och_count <= 0;
          conv2d_2_row_select <= 0;
          conv2d_2_prev_row_count <= 0;
          conv2d_2_prev_bat_count <= 0;
          conv2d_2_prev_och_count <= 0;
          conv2d_2_prev_row_select <= 0;
          conv2d_2_out_col_count <= 0;
          conv2d_2_out_row_count <= 0;
          conv2d_2_out_ram_select <= 0;
          conv2d_2_skip_read_filter <= 0;
          conv2d_2_skip_read_act <= 0;
          conv2d_2_skip_comp <= 0;
          conv2d_2_skip_write_out <= 1;
          if(cparam_conv2d_2_data_stationary == 0) begin
            control_conv2d_2 <= control_conv2d_2_3;
          end 
          if(cparam_conv2d_2_data_stationary == 1) begin
            control_conv2d_2 <= control_conv2d_2_8;
          end 
        end
        control_conv2d_2_3: begin
          control_conv2d_2 <= control_conv2d_2_4;
          if(conv2d_2_skip_read_filter) begin
            control_conv2d_2 <= control_conv2d_2_7;
          end 
        end
        control_conv2d_2_4: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_2 <= control_conv2d_2_5;
          end 
        end
        control_conv2d_2_5: begin
          if(_maxi_read_idle) begin
            control_conv2d_2 <= control_conv2d_2_6;
          end 
        end
        control_conv2d_2_6: begin
          control_conv2d_2 <= control_conv2d_2_7;
        end
        control_conv2d_2_7: begin
          if(cparam_conv2d_2_data_stationary == 0) begin
            control_conv2d_2 <= control_conv2d_2_8;
          end 
          if(cparam_conv2d_2_data_stationary == 1) begin
            control_conv2d_2 <= control_conv2d_2_20;
          end 
        end
        control_conv2d_2_8: begin
          control_conv2d_2 <= control_conv2d_2_9;
          if(conv2d_2_skip_read_act) begin
            control_conv2d_2 <= control_conv2d_2_19;
          end 
        end
        control_conv2d_2_9: begin
          control_conv2d_2 <= control_conv2d_2_10;
          if(conv2d_2_mux_dma_pad_mask_0 || !conv2d_2_mux_dma_flag_0) begin
            control_conv2d_2 <= control_conv2d_2_12;
          end 
        end
        control_conv2d_2_10: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_2 <= control_conv2d_2_11;
          end 
        end
        control_conv2d_2_11: begin
          if(_maxi_read_idle) begin
            control_conv2d_2 <= control_conv2d_2_12;
          end 
        end
        control_conv2d_2_12: begin
          control_conv2d_2 <= control_conv2d_2_13;
          if(conv2d_2_mux_dma_pad_mask_1 || !conv2d_2_mux_dma_flag_1) begin
            control_conv2d_2 <= control_conv2d_2_15;
          end 
        end
        control_conv2d_2_13: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_2 <= control_conv2d_2_14;
          end 
        end
        control_conv2d_2_14: begin
          if(_maxi_read_idle) begin
            control_conv2d_2 <= control_conv2d_2_15;
          end 
        end
        control_conv2d_2_15: begin
          control_conv2d_2 <= control_conv2d_2_16;
          if(conv2d_2_mux_dma_pad_mask_2 || !conv2d_2_mux_dma_flag_2) begin
            control_conv2d_2 <= control_conv2d_2_18;
          end 
        end
        control_conv2d_2_16: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_2 <= control_conv2d_2_17;
          end 
        end
        control_conv2d_2_17: begin
          if(_maxi_read_idle) begin
            control_conv2d_2 <= control_conv2d_2_18;
          end 
        end
        control_conv2d_2_18: begin
          control_conv2d_2 <= control_conv2d_2_19;
        end
        control_conv2d_2_19: begin
          if(cparam_conv2d_2_data_stationary == 0) begin
            control_conv2d_2 <= control_conv2d_2_20;
          end 
          if(cparam_conv2d_2_data_stationary == 1) begin
            control_conv2d_2 <= control_conv2d_2_3;
          end 
        end
        control_conv2d_2_20: begin
          if(_maxi_write_idle) begin
            control_conv2d_2 <= control_conv2d_2_21;
          end 
        end
        control_conv2d_2_21: begin
          if(conv2d_2_comp_fsm == 0) begin
            control_conv2d_2 <= control_conv2d_2_22;
          end 
        end
        control_conv2d_2_22: begin
          control_conv2d_2 <= control_conv2d_2_23;
          if(conv2d_2_skip_write_out) begin
            control_conv2d_2 <= control_conv2d_2_28;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_prev_och_count < cparam_conv2d_2_max_och_count)) begin
            control_conv2d_2 <= control_conv2d_2_28;
          end 
        end
        control_conv2d_2_23: begin
          if(conv2d_2_sync_comp_count >= conv2d_2_sync_out_count + cparam_conv2d_2_inc_sync_out) begin
            control_conv2d_2 <= control_conv2d_2_24;
          end 
        end
        control_conv2d_2_24: begin
          if(!conv2d_2_dma_out_mask_0) begin
            control_conv2d_2 <= control_conv2d_2_25;
          end 
          if(conv2d_2_dma_out_mask_0) begin
            control_conv2d_2 <= control_conv2d_2_26;
          end 
        end
        control_conv2d_2_25: begin
          if(_maxi_write_req_idle) begin
            control_conv2d_2 <= control_conv2d_2_26;
          end 
        end
        control_conv2d_2_26: begin
          control_conv2d_2 <= control_conv2d_2_27;
        end
        control_conv2d_2_27: begin
          conv2d_2_write_count <= conv2d_2_write_count + 1;
          if(conv2d_2_out_ram_select == 0) begin
            conv2d_2_out_laddr_offset <= conv2d_2_out_laddr_offset + conv2d_2_next_out_write_size;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && !cparam_conv2d_2_keep_filter) begin
            conv2d_2_out_base_offset_col <= conv2d_2_out_base_offset_col + cparam_conv2d_2_out_col_step;
            conv2d_2_out_col_count <= conv2d_2_out_col_count + 1;
          end 
          conv2d_2_out_ram_select <= conv2d_2_out_ram_select + 1;
          if(conv2d_2_out_ram_select == 0) begin
            conv2d_2_out_ram_select <= 0;
          end 
          conv2d_2_sync_out_count <= conv2d_2_sync_out_count + cparam_conv2d_2_inc_sync_out;
          if((cparam_conv2d_2_data_stationary == 0) && !cparam_conv2d_2_keep_filter && (conv2d_2_write_count >= cparam_conv2d_2_out_num_col - 1) || (cparam_conv2d_2_data_stationary == 0) && cparam_conv2d_2_keep_filter || (cparam_conv2d_2_data_stationary == 1)) begin
            conv2d_2_sync_out_count <= conv2d_2_sync_out_count + (cparam_conv2d_2_inc_sync_out + cparam_conv2d_2_inc_sync_out_res);
          end 
          if((cparam_conv2d_2_data_stationary == 0) && !cparam_conv2d_2_keep_filter) begin
            control_conv2d_2 <= control_conv2d_2_22;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && !cparam_conv2d_2_keep_filter && (conv2d_2_write_count >= cparam_conv2d_2_out_num_col - 1) || (cparam_conv2d_2_data_stationary == 0) && cparam_conv2d_2_keep_filter || (cparam_conv2d_2_data_stationary == 1)) begin
            control_conv2d_2 <= control_conv2d_2_28;
          end 
        end
        control_conv2d_2_28: begin
          if(conv2d_2_update_filter) begin
            conv2d_2_filter_base_offset <= conv2d_2_filter_base_offset + cparam_conv2d_2_filter_base_step;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)) begin
            conv2d_2_filter_base_offset <= 0;
          end 
          if(conv2d_2_update_filter) begin
            conv2d_2_och_count <= conv2d_2_och_count + cparam_conv2d_2_och_count_step;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)) begin
            conv2d_2_och_count <= 0;
          end 
          if(conv2d_2_update_filter) begin
            conv2d_2_filter_page_comp_offset <= conv2d_2_filter_page_comp_offset + cparam_conv2d_2_filter_read_step;
            conv2d_2_filter_page_dma_offset <= conv2d_2_filter_page_dma_offset + cparam_conv2d_2_filter_read_step;
          end 
          if(conv2d_2_update_filter && (conv2d_2_filter_page_comp_offset + cparam_conv2d_2_filter_read_step + cparam_conv2d_2_filter_read_step > 128)) begin
            conv2d_2_filter_page_comp_offset <= 0;
            conv2d_2_filter_page_dma_offset <= 0;
          end 
          if(conv2d_2_update_act) begin
            conv2d_2_act_base_offset_row <= conv2d_2_act_base_offset_row + cparam_conv2d_2_act_row_step;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)) begin
            conv2d_2_act_base_offset_row <= 0;
            conv2d_2_act_base_offset_bat <= conv2d_2_act_base_offset_bat + cparam_conv2d_2_act_bat_step;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count)) begin
            conv2d_2_act_base_offset_bat <= 0;
          end 
          if(!conv2d_2_update_act) begin
            conv2d_2_dma_flag_0 <= 0;
          end 
          if(conv2d_2_update_act) begin
            conv2d_2_dma_flag_0 <= cparam_conv2d_2_dma_flag_conds_0;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)) begin
            conv2d_2_dma_flag_0 <= 1;
          end 
          if(!conv2d_2_update_act) begin
            conv2d_2_dma_flag_1 <= 0;
          end 
          if(conv2d_2_update_act) begin
            conv2d_2_dma_flag_1 <= cparam_conv2d_2_dma_flag_conds_1;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)) begin
            conv2d_2_dma_flag_1 <= 1;
          end 
          if(!conv2d_2_update_act) begin
            conv2d_2_dma_flag_2 <= 0;
          end 
          if(conv2d_2_update_act) begin
            conv2d_2_dma_flag_2 <= cparam_conv2d_2_dma_flag_conds_2;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)) begin
            conv2d_2_dma_flag_2 <= 1;
          end 
          if(conv2d_2_update_act) begin
            conv2d_2_row_count <= conv2d_2_row_count + cparam_conv2d_2_stride_row_par_row;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)) begin
            conv2d_2_row_count <= 0;
            conv2d_2_bat_count <= conv2d_2_bat_count + 1;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count)) begin
            conv2d_2_bat_count <= 0;
          end 
          if(conv2d_2_update_act && (cparam_conv2d_2_stride_row_par_row < 3)) begin
            conv2d_2_row_select <= conv2d_2_row_select + cparam_conv2d_2_stride_row_par_row;
            conv2d_2_prev_row_select <= conv2d_2_row_select;
          end 
          if(conv2d_2_update_act && (cparam_conv2d_2_stride_row_par_row < 3) && (conv2d_2_row_select + cparam_conv2d_2_stride_row_par_row >= 3)) begin
            conv2d_2_row_select <= conv2d_2_row_select - (3 - cparam_conv2d_2_stride_row_par_row);
            conv2d_2_prev_row_select <= conv2d_2_row_select;
          end 
          if(conv2d_2_update_act && !(cparam_conv2d_2_stride_row_par_row < 3)) begin
            conv2d_2_row_select <= 0;
            conv2d_2_prev_row_select <= 0;
          end 
          if(conv2d_2_update_act && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count)) begin
            conv2d_2_row_select <= 0;
            conv2d_2_prev_row_select <= 0;
          end 
          if(conv2d_2_update_act && conv2d_2_mux_next_dma_flag_0) begin
            conv2d_2_act_page_comp_offset_0 <= conv2d_2_act_page_comp_offset_0 + cparam_conv2d_2_act_read_step;
            conv2d_2_act_page_dma_offset_0 <= conv2d_2_act_page_dma_offset_0 + cparam_conv2d_2_act_read_step;
          end 
          if(conv2d_2_update_act && conv2d_2_mux_next_dma_flag_0 && (conv2d_2_act_page_comp_offset_0 + cparam_conv2d_2_act_read_step + cparam_conv2d_2_act_read_step > 128)) begin
            conv2d_2_act_page_comp_offset_0 <= 0;
            conv2d_2_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) && cparam_conv2d_2_keep_input) begin
            conv2d_2_act_page_comp_offset_0 <= 0;
            conv2d_2_act_page_dma_offset_0 <= 0;
          end 
          if(conv2d_2_update_act && conv2d_2_mux_next_dma_flag_1) begin
            conv2d_2_act_page_comp_offset_1 <= conv2d_2_act_page_comp_offset_1 + cparam_conv2d_2_act_read_step;
            conv2d_2_act_page_dma_offset_1 <= conv2d_2_act_page_dma_offset_1 + cparam_conv2d_2_act_read_step;
          end 
          if(conv2d_2_update_act && conv2d_2_mux_next_dma_flag_1 && (conv2d_2_act_page_comp_offset_1 + cparam_conv2d_2_act_read_step + cparam_conv2d_2_act_read_step > 128)) begin
            conv2d_2_act_page_comp_offset_1 <= 0;
            conv2d_2_act_page_dma_offset_1 <= 0;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) && cparam_conv2d_2_keep_input) begin
            conv2d_2_act_page_comp_offset_1 <= 0;
            conv2d_2_act_page_dma_offset_1 <= 0;
          end 
          if(conv2d_2_update_act && conv2d_2_mux_next_dma_flag_2) begin
            conv2d_2_act_page_comp_offset_2 <= conv2d_2_act_page_comp_offset_2 + cparam_conv2d_2_act_read_step;
            conv2d_2_act_page_dma_offset_2 <= conv2d_2_act_page_dma_offset_2 + cparam_conv2d_2_act_read_step;
          end 
          if(conv2d_2_update_act && conv2d_2_mux_next_dma_flag_2 && (conv2d_2_act_page_comp_offset_2 + cparam_conv2d_2_act_read_step + cparam_conv2d_2_act_read_step > 128)) begin
            conv2d_2_act_page_comp_offset_2 <= 0;
            conv2d_2_act_page_dma_offset_2 <= 0;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) && cparam_conv2d_2_keep_input) begin
            conv2d_2_act_page_comp_offset_2 <= 0;
            conv2d_2_act_page_dma_offset_2 <= 0;
          end 
          conv2d_2_next_out_write_size <= (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)? cparam_conv2d_2_out_write_size_res : cparam_conv2d_2_out_write_size;
          if(!conv2d_2_skip_write_out) begin
            conv2d_2_write_count <= 0;
            conv2d_2_out_laddr_offset <= 0;
            conv2d_2_out_ram_select <= 0;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && !conv2d_2_skip_write_out) begin
            conv2d_2_out_base_offset_col <= 0;
            conv2d_2_out_base_offset_row <= conv2d_2_out_base_offset_row + cparam_conv2d_2_out_row_step;
            conv2d_2_out_col_count <= 0;
            conv2d_2_out_row_count <= conv2d_2_out_row_count + 1;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && !conv2d_2_skip_write_out && (conv2d_2_prev_row_count >= cparam_conv2d_2_max_row_count)) begin
            conv2d_2_out_base_offset_row <= 0;
            conv2d_2_out_base_offset_bat <= conv2d_2_out_base_offset_bat + cparam_conv2d_2_out_bat_step;
            conv2d_2_out_row_count <= 0;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && !conv2d_2_skip_write_out && (conv2d_2_prev_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_prev_bat_count >= cparam_conv2d_2_max_bat_count)) begin
            conv2d_2_out_base_offset_bat <= 0;
            conv2d_2_out_base_offset_och <= conv2d_2_out_base_offset_och + cparam_conv2d_2_out_och_step;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_prev_och_count >= cparam_conv2d_2_max_och_count) && !conv2d_2_skip_write_out) begin
            conv2d_2_out_base_offset_row <= conv2d_2_out_base_offset_row + cparam_conv2d_2_out_row_step;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && !conv2d_2_out_page) begin
            conv2d_2_out_page_comp_offset <= 64;
            conv2d_2_out_page_dma_offset <= 0;
            conv2d_2_out_page <= 1;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && conv2d_2_out_page) begin
            conv2d_2_out_page_comp_offset <= 0;
            conv2d_2_out_page_dma_offset <= 64;
            conv2d_2_out_page <= 0;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count) && !conv2d_2_out_page) begin
            conv2d_2_out_page_comp_offset <= 64;
            conv2d_2_out_page_dma_offset <= 0;
            conv2d_2_out_page <= 1;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count) && conv2d_2_out_page) begin
            conv2d_2_out_page_comp_offset <= 0;
            conv2d_2_out_page_dma_offset <= 64;
            conv2d_2_out_page <= 0;
          end 
          conv2d_2_prev_row_count <= conv2d_2_row_count;
          conv2d_2_prev_bat_count <= conv2d_2_bat_count;
          conv2d_2_prev_och_count <= conv2d_2_och_count;
          if((conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)) begin
            conv2d_2_skip_read_filter <= 1;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && cparam_conv2d_2_keep_filter) begin
            conv2d_2_skip_read_filter <= 1;
          end 
          if((conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)) begin
            conv2d_2_skip_read_act <= 1;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) && cparam_conv2d_2_keep_input) begin
            conv2d_2_skip_read_act <= 1;
          end 
          if((conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)) begin
            conv2d_2_skip_comp <= 1;
          end 
          if(conv2d_2_skip_write_out && (conv2d_2_prev_row_count == 0) && (conv2d_2_prev_bat_count == 0) && (conv2d_2_prev_och_count == 0)) begin
            conv2d_2_skip_write_out <= 0;
          end 
          if(cparam_conv2d_2_data_stationary == 0) begin
            control_conv2d_2 <= control_conv2d_2_8;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && (conv2d_2_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_bat_count >= cparam_conv2d_2_max_bat_count)) begin
            control_conv2d_2 <= control_conv2d_2_3;
          end 
          if(cparam_conv2d_2_data_stationary == 1) begin
            control_conv2d_2 <= control_conv2d_2_3;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)) begin
            control_conv2d_2 <= control_conv2d_2_8;
          end 
          if(!conv2d_2_skip_write_out && (conv2d_2_prev_och_count >= cparam_conv2d_2_max_och_count) && (conv2d_2_prev_row_count >= cparam_conv2d_2_max_row_count) && (conv2d_2_prev_bat_count >= cparam_conv2d_2_max_bat_count)) begin
            control_conv2d_2 <= control_conv2d_2_29;
          end 
        end
        control_conv2d_2_29: begin
          if(_maxi_write_idle && (outstanding_wcount_0 == 0)) begin
            control_conv2d_2 <= control_conv2d_2_30;
          end 
        end
        control_conv2d_2_30: begin
          if(main_fsm == 11) begin
            _control_conv2d_2_called <= 0;
          end 
          if(main_fsm == 11) begin
            control_conv2d_2 <= control_conv2d_2_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
      _maxi_read_cont <= 0;
    end else begin
      case(_maxi_read_req_fsm)
        _maxi_read_req_fsm_init: begin
          if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_1;
          end 
        end
        _maxi_read_req_fsm_1: begin
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_cont <= 1;
          end 
          if((maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
            _maxi_read_cont <= 0;
          end 
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_data_fsm_1 = 1;
  localparam _maxi_read_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
    end else begin
      case(_maxi_read_data_fsm)
        _maxi_read_data_fsm_init: begin
          if(_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(_maxi_read_data_idle && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
        end
        _maxi_read_data_fsm_1: begin
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
        end
        _maxi_read_data_fsm_2: begin
          if(maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(maxi_rvalid && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_0_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_0 <= write_burst_fsm_0_init;
      write_burst_addr_49 <= 0;
      write_burst_stride_50 <= 0;
      write_burst_length_51 <= 0;
      write_burst_done_52 <= 0;
    end else begin
      case(write_burst_fsm_0)
        write_burst_fsm_0_init: begin
          write_burst_addr_49 <= _maxi_read_local_addr_buf;
          write_burst_stride_50 <= _maxi_read_local_stride_buf;
          write_burst_length_51 <= _maxi_read_local_size_buf;
          write_burst_done_52 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_1;
          end 
        end
        write_burst_fsm_0_1: begin
          if(write_burst_block_ram_wvalid_47) begin
            write_burst_addr_49 <= write_burst_addr_49 + write_burst_stride_50;
            write_burst_length_51 <= write_burst_length_51 - 1;
            write_burst_done_52 <= 0;
          end 
          if(write_burst_block_ram_wvalid_47 && (write_burst_length_51 <= 1)) begin
            write_burst_done_52 <= 1;
          end 
          if(write_burst_block_ram_wvalid_47 && 0) begin
            write_burst_done_52 <= 1;
          end 
          if(write_burst_block_ram_wvalid_47 && (write_burst_length_51 <= 1)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(write_burst_block_ram_wvalid_47 && 0) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(write_burst_block_ram_wquit_48) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_1_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_1 <= write_burst_fsm_1_init;
      write_burst_addr_55 <= 0;
      write_burst_stride_56 <= 0;
      write_burst_length_57 <= 0;
      write_burst_done_58 <= 0;
    end else begin
      case(write_burst_fsm_1)
        write_burst_fsm_1_init: begin
          write_burst_addr_55 <= _maxi_read_local_addr_buf;
          write_burst_stride_56 <= _maxi_read_local_stride_buf;
          write_burst_length_57 <= _maxi_read_local_size_buf;
          write_burst_done_58 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_1 <= write_burst_fsm_1_1;
          end 
        end
        write_burst_fsm_1_1: begin
          if(write_burst_block_ram_wvalid_53) begin
            write_burst_addr_55 <= write_burst_addr_55 + write_burst_stride_56;
            write_burst_length_57 <= write_burst_length_57 - 1;
            write_burst_done_58 <= 0;
          end 
          if(write_burst_block_ram_wvalid_53 && (write_burst_length_57 <= 1)) begin
            write_burst_done_58 <= 1;
          end 
          if(write_burst_block_ram_wvalid_53 && 0) begin
            write_burst_done_58 <= 1;
          end 
          if(write_burst_block_ram_wvalid_53 && (write_burst_length_57 <= 1)) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
          if(write_burst_block_ram_wvalid_53 && 0) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
          if(write_burst_block_ram_wquit_54) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_2_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_2 <= write_burst_fsm_2_init;
      write_burst_addr_61 <= 0;
      write_burst_stride_62 <= 0;
      write_burst_length_63 <= 0;
      write_burst_done_64 <= 0;
    end else begin
      case(write_burst_fsm_2)
        write_burst_fsm_2_init: begin
          write_burst_addr_61 <= _maxi_read_local_addr_buf;
          write_burst_stride_62 <= _maxi_read_local_stride_buf;
          write_burst_length_63 <= _maxi_read_local_size_buf;
          write_burst_done_64 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_1;
          end 
        end
        write_burst_fsm_2_1: begin
          if(write_burst_block_ram_wvalid_59) begin
            write_burst_addr_61 <= write_burst_addr_61 + write_burst_stride_62;
            write_burst_length_63 <= write_burst_length_63 - 1;
            write_burst_done_64 <= 0;
          end 
          if(write_burst_block_ram_wvalid_59 && (write_burst_length_63 <= 1)) begin
            write_burst_done_64 <= 1;
          end 
          if(write_burst_block_ram_wvalid_59 && 0) begin
            write_burst_done_64 <= 1;
          end 
          if(write_burst_block_ram_wvalid_59 && (write_burst_length_63 <= 1)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(write_burst_block_ram_wvalid_59 && 0) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(write_burst_block_ram_wquit_60) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_3_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_3 <= write_burst_fsm_3_init;
      write_burst_addr_67 <= 0;
      write_burst_stride_68 <= 0;
      write_burst_length_69 <= 0;
      write_burst_done_70 <= 0;
    end else begin
      case(write_burst_fsm_3)
        write_burst_fsm_3_init: begin
          write_burst_addr_67 <= _maxi_read_local_addr_buf;
          write_burst_stride_68 <= _maxi_read_local_stride_buf;
          write_burst_length_69 <= _maxi_read_local_size_buf;
          write_burst_done_70 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_1;
          end 
        end
        write_burst_fsm_3_1: begin
          if(write_burst_block_ram_wvalid_65) begin
            write_burst_addr_67 <= write_burst_addr_67 + write_burst_stride_68;
            write_burst_length_69 <= write_burst_length_69 - 1;
            write_burst_done_70 <= 0;
          end 
          if(write_burst_block_ram_wvalid_65 && (write_burst_length_69 <= 1)) begin
            write_burst_done_70 <= 1;
          end 
          if(write_burst_block_ram_wvalid_65 && 0) begin
            write_burst_done_70 <= 1;
          end 
          if(write_burst_block_ram_wvalid_65 && (write_burst_length_69 <= 1)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(write_burst_block_ram_wvalid_65 && 0) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(write_burst_block_ram_wquit_66) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_4_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_4 <= write_burst_fsm_4_init;
      write_burst_addr_73 <= 0;
      write_burst_stride_74 <= 0;
      write_burst_length_75 <= 0;
      write_burst_done_76 <= 0;
    end else begin
      case(write_burst_fsm_4)
        write_burst_fsm_4_init: begin
          write_burst_addr_73 <= _maxi_read_local_addr_buf;
          write_burst_stride_74 <= _maxi_read_local_stride_buf;
          write_burst_length_75 <= _maxi_read_local_size_buf;
          write_burst_done_76 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_4 <= write_burst_fsm_4_1;
          end 
        end
        write_burst_fsm_4_1: begin
          if(write_burst_block_ram_wvalid_71) begin
            write_burst_addr_73 <= write_burst_addr_73 + write_burst_stride_74;
            write_burst_length_75 <= write_burst_length_75 - 1;
            write_burst_done_76 <= 0;
          end 
          if(write_burst_block_ram_wvalid_71 && (write_burst_length_75 <= 1)) begin
            write_burst_done_76 <= 1;
          end 
          if(write_burst_block_ram_wvalid_71 && 0) begin
            write_burst_done_76 <= 1;
          end 
          if(write_burst_block_ram_wvalid_71 && (write_burst_length_75 <= 1)) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
          if(write_burst_block_ram_wvalid_71 && 0) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
          if(write_burst_block_ram_wquit_72) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_5_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_5 <= write_burst_fsm_5_init;
      write_burst_addr_79 <= 0;
      write_burst_stride_80 <= 0;
      write_burst_length_81 <= 0;
      write_burst_done_82 <= 0;
    end else begin
      case(write_burst_fsm_5)
        write_burst_fsm_5_init: begin
          write_burst_addr_79 <= _maxi_read_local_addr_buf;
          write_burst_stride_80 <= _maxi_read_local_stride_buf;
          write_burst_length_81 <= _maxi_read_local_size_buf;
          write_burst_done_82 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_5 <= write_burst_fsm_5_1;
          end 
        end
        write_burst_fsm_5_1: begin
          if(write_burst_block_ram_wvalid_77) begin
            write_burst_addr_79 <= write_burst_addr_79 + write_burst_stride_80;
            write_burst_length_81 <= write_burst_length_81 - 1;
            write_burst_done_82 <= 0;
          end 
          if(write_burst_block_ram_wvalid_77 && (write_burst_length_81 <= 1)) begin
            write_burst_done_82 <= 1;
          end 
          if(write_burst_block_ram_wvalid_77 && 0) begin
            write_burst_done_82 <= 1;
          end 
          if(write_burst_block_ram_wvalid_77 && (write_burst_length_81 <= 1)) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
          if(write_burst_block_ram_wvalid_77 && 0) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
          if(write_burst_block_ram_wquit_78) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_6_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_6 <= write_burst_fsm_6_init;
      write_burst_addr_85 <= 0;
      write_burst_stride_86 <= 0;
      write_burst_length_87 <= 0;
      write_burst_done_88 <= 0;
    end else begin
      case(write_burst_fsm_6)
        write_burst_fsm_6_init: begin
          write_burst_addr_85 <= _maxi_read_local_addr_buf;
          write_burst_stride_86 <= _maxi_read_local_stride_buf;
          write_burst_length_87 <= _maxi_read_local_size_buf;
          write_burst_done_88 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_6 <= write_burst_fsm_6_1;
          end 
        end
        write_burst_fsm_6_1: begin
          if(write_burst_block_ram_wvalid_83) begin
            write_burst_addr_85 <= write_burst_addr_85 + write_burst_stride_86;
            write_burst_length_87 <= write_burst_length_87 - 1;
            write_burst_done_88 <= 0;
          end 
          if(write_burst_block_ram_wvalid_83 && (write_burst_length_87 <= 1)) begin
            write_burst_done_88 <= 1;
          end 
          if(write_burst_block_ram_wvalid_83 && 0) begin
            write_burst_done_88 <= 1;
          end 
          if(write_burst_block_ram_wvalid_83 && (write_burst_length_87 <= 1)) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
          if(write_burst_block_ram_wvalid_83 && 0) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
          if(write_burst_block_ram_wquit_84) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_7_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_7 <= write_burst_fsm_7_init;
      write_burst_addr_91 <= 0;
      write_burst_stride_92 <= 0;
      write_burst_length_93 <= 0;
      write_burst_done_94 <= 0;
    end else begin
      case(write_burst_fsm_7)
        write_burst_fsm_7_init: begin
          write_burst_addr_91 <= _maxi_read_local_addr_buf;
          write_burst_stride_92 <= _maxi_read_local_stride_buf;
          write_burst_length_93 <= _maxi_read_local_size_buf;
          write_burst_done_94 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_7 <= write_burst_fsm_7_1;
          end 
        end
        write_burst_fsm_7_1: begin
          if(write_burst_block_ram_wvalid_89) begin
            write_burst_addr_91 <= write_burst_addr_91 + write_burst_stride_92;
            write_burst_length_93 <= write_burst_length_93 - 1;
            write_burst_done_94 <= 0;
          end 
          if(write_burst_block_ram_wvalid_89 && (write_burst_length_93 <= 1)) begin
            write_burst_done_94 <= 1;
          end 
          if(write_burst_block_ram_wvalid_89 && 0) begin
            write_burst_done_94 <= 1;
          end 
          if(write_burst_block_ram_wvalid_89 && (write_burst_length_93 <= 1)) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
          if(write_burst_block_ram_wvalid_89 && 0) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
          if(write_burst_block_ram_wquit_90) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_8_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_8 <= write_burst_fsm_8_init;
      write_burst_addr_97 <= 0;
      write_burst_stride_98 <= 0;
      write_burst_length_99 <= 0;
      write_burst_done_100 <= 0;
    end else begin
      case(write_burst_fsm_8)
        write_burst_fsm_8_init: begin
          write_burst_addr_97 <= _maxi_read_local_addr_buf;
          write_burst_stride_98 <= _maxi_read_local_stride_buf;
          write_burst_length_99 <= _maxi_read_local_size_buf;
          write_burst_done_100 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_8 <= write_burst_fsm_8_1;
          end 
        end
        write_burst_fsm_8_1: begin
          if(write_burst_block_ram_wvalid_95) begin
            write_burst_addr_97 <= write_burst_addr_97 + write_burst_stride_98;
            write_burst_length_99 <= write_burst_length_99 - 1;
            write_burst_done_100 <= 0;
          end 
          if(write_burst_block_ram_wvalid_95 && (write_burst_length_99 <= 1)) begin
            write_burst_done_100 <= 1;
          end 
          if(write_burst_block_ram_wvalid_95 && 0) begin
            write_burst_done_100 <= 1;
          end 
          if(write_burst_block_ram_wvalid_95 && (write_burst_length_99 <= 1)) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
          if(write_burst_block_ram_wvalid_95 && 0) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
          if(write_burst_block_ram_wquit_96) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_9_1 = 1;
  localparam write_burst_block_fsm_9_2 = 2;
  localparam write_burst_block_fsm_9_3 = 3;
  localparam write_burst_block_fsm_9_4 = 4;
  localparam write_burst_block_fsm_9_5 = 5;
  localparam write_burst_block_fsm_9_6 = 6;
  localparam write_burst_block_fsm_9_7 = 7;
  localparam write_burst_block_fsm_9_8 = 8;
  localparam write_burst_block_fsm_9_9 = 9;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
      write_burst_block_length_101 <= 0;
      write_burst_block_blocksize_102 <= 0;
      write_burst_block_done_103 <= 0;
      write_burst_block_count_104 <= 0;
    end else begin
      case(write_burst_block_fsm_9)
        write_burst_block_fsm_9_init: begin
          write_burst_block_length_101 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_102 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_103 <= 0;
          write_burst_block_count_104 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_1;
          end 
        end
        write_burst_block_fsm_9_1: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_2;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_2: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_3;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_3: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_4;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_4: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_5;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_5: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_6;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_6: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_7;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_7: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_8;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_8: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_9;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
        write_burst_block_fsm_9_9: begin
          if(maxi_rvalid) begin
            write_burst_block_length_101 <= write_burst_block_length_101 - 1;
            write_burst_block_done_103 <= 0;
            write_burst_block_count_104 <= write_burst_block_count_104 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_103 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_count_104 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_104 == write_burst_block_blocksize_102 - 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_1;
          end 
          if(maxi_rvalid && (write_burst_block_length_101 <= 1)) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
          if(0) begin
            write_burst_block_fsm_9 <= write_burst_block_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_10_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_10 <= write_burst_fsm_10_init;
      write_burst_addr_109 <= 0;
      write_burst_stride_110 <= 0;
      write_burst_length_111 <= 0;
      write_burst_done_112 <= 0;
    end else begin
      case(write_burst_fsm_10)
        write_burst_fsm_10_init: begin
          write_burst_addr_109 <= _maxi_read_local_addr_buf;
          write_burst_stride_110 <= _maxi_read_local_stride_buf;
          write_burst_length_111 <= _maxi_read_local_size_buf;
          write_burst_done_112 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_10 <= write_burst_fsm_10_1;
          end 
        end
        write_burst_fsm_10_1: begin
          if(write_burst_block_ram_wvalid_107) begin
            write_burst_addr_109 <= write_burst_addr_109 + write_burst_stride_110;
            write_burst_length_111 <= write_burst_length_111 - 1;
            write_burst_done_112 <= 0;
          end 
          if(write_burst_block_ram_wvalid_107 && (write_burst_length_111 <= 1)) begin
            write_burst_done_112 <= 1;
          end 
          if(write_burst_block_ram_wvalid_107 && 0) begin
            write_burst_done_112 <= 1;
          end 
          if(write_burst_block_ram_wvalid_107 && (write_burst_length_111 <= 1)) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
          if(write_burst_block_ram_wvalid_107 && 0) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
          if(write_burst_block_ram_wquit_108) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_11_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_11 <= write_burst_fsm_11_init;
      write_burst_addr_115 <= 0;
      write_burst_stride_116 <= 0;
      write_burst_length_117 <= 0;
      write_burst_done_118 <= 0;
    end else begin
      case(write_burst_fsm_11)
        write_burst_fsm_11_init: begin
          write_burst_addr_115 <= _maxi_read_local_addr_buf;
          write_burst_stride_116 <= _maxi_read_local_stride_buf;
          write_burst_length_117 <= _maxi_read_local_size_buf;
          write_burst_done_118 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_11 <= write_burst_fsm_11_1;
          end 
        end
        write_burst_fsm_11_1: begin
          if(write_burst_block_ram_wvalid_113) begin
            write_burst_addr_115 <= write_burst_addr_115 + write_burst_stride_116;
            write_burst_length_117 <= write_burst_length_117 - 1;
            write_burst_done_118 <= 0;
          end 
          if(write_burst_block_ram_wvalid_113 && (write_burst_length_117 <= 1)) begin
            write_burst_done_118 <= 1;
          end 
          if(write_burst_block_ram_wvalid_113 && 0) begin
            write_burst_done_118 <= 1;
          end 
          if(write_burst_block_ram_wvalid_113 && (write_burst_length_117 <= 1)) begin
            write_burst_fsm_11 <= write_burst_fsm_11_init;
          end 
          if(write_burst_block_ram_wvalid_113 && 0) begin
            write_burst_fsm_11 <= write_burst_fsm_11_init;
          end 
          if(write_burst_block_ram_wquit_114) begin
            write_burst_fsm_11 <= write_burst_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_12_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_12 <= write_burst_fsm_12_init;
      write_burst_addr_121 <= 0;
      write_burst_stride_122 <= 0;
      write_burst_length_123 <= 0;
      write_burst_done_124 <= 0;
    end else begin
      case(write_burst_fsm_12)
        write_burst_fsm_12_init: begin
          write_burst_addr_121 <= _maxi_read_local_addr_buf;
          write_burst_stride_122 <= _maxi_read_local_stride_buf;
          write_burst_length_123 <= _maxi_read_local_size_buf;
          write_burst_done_124 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_12 <= write_burst_fsm_12_1;
          end 
        end
        write_burst_fsm_12_1: begin
          if(write_burst_block_ram_wvalid_119) begin
            write_burst_addr_121 <= write_burst_addr_121 + write_burst_stride_122;
            write_burst_length_123 <= write_burst_length_123 - 1;
            write_burst_done_124 <= 0;
          end 
          if(write_burst_block_ram_wvalid_119 && (write_burst_length_123 <= 1)) begin
            write_burst_done_124 <= 1;
          end 
          if(write_burst_block_ram_wvalid_119 && 0) begin
            write_burst_done_124 <= 1;
          end 
          if(write_burst_block_ram_wvalid_119 && (write_burst_length_123 <= 1)) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
          if(write_burst_block_ram_wvalid_119 && 0) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
          if(write_burst_block_ram_wquit_120) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_13_1 = 1;
  localparam write_burst_block_fsm_13_2 = 2;
  localparam write_burst_block_fsm_13_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
      write_burst_block_length_125 <= 0;
      write_burst_block_blocksize_126 <= 0;
      write_burst_block_done_127 <= 0;
      write_burst_block_count_128 <= 0;
    end else begin
      case(write_burst_block_fsm_13)
        write_burst_block_fsm_13_init: begin
          write_burst_block_length_125 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_126 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_127 <= 0;
          write_burst_block_count_128 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_1;
          end 
        end
        write_burst_block_fsm_13_1: begin
          if(maxi_rvalid) begin
            write_burst_block_length_125 <= write_burst_block_length_125 - 1;
            write_burst_block_done_127 <= 0;
            write_burst_block_count_128 <= write_burst_block_count_128 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_125 <= 1)) begin
            write_burst_block_done_127 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_127 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_128 == write_burst_block_blocksize_126 - 1)) begin
            write_burst_block_count_128 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_128 == write_burst_block_blocksize_126 - 1)) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_2;
          end 
          if(maxi_rvalid && (write_burst_block_length_125 <= 1)) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
          if(0) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
        end
        write_burst_block_fsm_13_2: begin
          if(maxi_rvalid) begin
            write_burst_block_length_125 <= write_burst_block_length_125 - 1;
            write_burst_block_done_127 <= 0;
            write_burst_block_count_128 <= write_burst_block_count_128 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_125 <= 1)) begin
            write_burst_block_done_127 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_127 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_128 == write_burst_block_blocksize_126 - 1)) begin
            write_burst_block_count_128 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_128 == write_burst_block_blocksize_126 - 1)) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_3;
          end 
          if(maxi_rvalid && (write_burst_block_length_125 <= 1)) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
          if(0) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
        end
        write_burst_block_fsm_13_3: begin
          if(maxi_rvalid) begin
            write_burst_block_length_125 <= write_burst_block_length_125 - 1;
            write_burst_block_done_127 <= 0;
            write_burst_block_count_128 <= write_burst_block_count_128 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_125 <= 1)) begin
            write_burst_block_done_127 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_127 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_128 == write_burst_block_blocksize_126 - 1)) begin
            write_burst_block_count_128 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_128 == write_burst_block_blocksize_126 - 1)) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_1;
          end 
          if(maxi_rvalid && (write_burst_block_length_125 <= 1)) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
          if(0) begin
            write_burst_block_fsm_13 <= write_burst_block_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_14_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_14 <= write_burst_fsm_14_init;
      write_burst_addr_133 <= 0;
      write_burst_stride_134 <= 0;
      write_burst_length_135 <= 0;
      write_burst_done_136 <= 0;
    end else begin
      case(write_burst_fsm_14)
        write_burst_fsm_14_init: begin
          write_burst_addr_133 <= _maxi_read_local_addr_buf;
          write_burst_stride_134 <= _maxi_read_local_stride_buf;
          write_burst_length_135 <= _maxi_read_local_size_buf;
          write_burst_done_136 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_14 <= write_burst_fsm_14_1;
          end 
        end
        write_burst_fsm_14_1: begin
          if(write_burst_block_ram_wvalid_131) begin
            write_burst_addr_133 <= write_burst_addr_133 + write_burst_stride_134;
            write_burst_length_135 <= write_burst_length_135 - 1;
            write_burst_done_136 <= 0;
          end 
          if(write_burst_block_ram_wvalid_131 && (write_burst_length_135 <= 1)) begin
            write_burst_done_136 <= 1;
          end 
          if(write_burst_block_ram_wvalid_131 && 0) begin
            write_burst_done_136 <= 1;
          end 
          if(write_burst_block_ram_wvalid_131 && (write_burst_length_135 <= 1)) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
          if(write_burst_block_ram_wvalid_131 && 0) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
          if(write_burst_block_ram_wquit_132) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_15_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_15 <= write_burst_fsm_15_init;
      write_burst_addr_139 <= 0;
      write_burst_stride_140 <= 0;
      write_burst_length_141 <= 0;
      write_burst_done_142 <= 0;
    end else begin
      case(write_burst_fsm_15)
        write_burst_fsm_15_init: begin
          write_burst_addr_139 <= _maxi_read_local_addr_buf;
          write_burst_stride_140 <= _maxi_read_local_stride_buf;
          write_burst_length_141 <= _maxi_read_local_size_buf;
          write_burst_done_142 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_15 <= write_burst_fsm_15_1;
          end 
        end
        write_burst_fsm_15_1: begin
          if(write_burst_block_ram_wvalid_137) begin
            write_burst_addr_139 <= write_burst_addr_139 + write_burst_stride_140;
            write_burst_length_141 <= write_burst_length_141 - 1;
            write_burst_done_142 <= 0;
          end 
          if(write_burst_block_ram_wvalid_137 && (write_burst_length_141 <= 1)) begin
            write_burst_done_142 <= 1;
          end 
          if(write_burst_block_ram_wvalid_137 && 0) begin
            write_burst_done_142 <= 1;
          end 
          if(write_burst_block_ram_wvalid_137 && (write_burst_length_141 <= 1)) begin
            write_burst_fsm_15 <= write_burst_fsm_15_init;
          end 
          if(write_burst_block_ram_wvalid_137 && 0) begin
            write_burst_fsm_15 <= write_burst_fsm_15_init;
          end 
          if(write_burst_block_ram_wquit_138) begin
            write_burst_fsm_15 <= write_burst_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_16_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_16 <= write_burst_fsm_16_init;
      write_burst_addr_145 <= 0;
      write_burst_stride_146 <= 0;
      write_burst_length_147 <= 0;
      write_burst_done_148 <= 0;
    end else begin
      case(write_burst_fsm_16)
        write_burst_fsm_16_init: begin
          write_burst_addr_145 <= _maxi_read_local_addr_buf;
          write_burst_stride_146 <= _maxi_read_local_stride_buf;
          write_burst_length_147 <= _maxi_read_local_size_buf;
          write_burst_done_148 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_16 <= write_burst_fsm_16_1;
          end 
        end
        write_burst_fsm_16_1: begin
          if(write_burst_block_ram_wvalid_143) begin
            write_burst_addr_145 <= write_burst_addr_145 + write_burst_stride_146;
            write_burst_length_147 <= write_burst_length_147 - 1;
            write_burst_done_148 <= 0;
          end 
          if(write_burst_block_ram_wvalid_143 && (write_burst_length_147 <= 1)) begin
            write_burst_done_148 <= 1;
          end 
          if(write_burst_block_ram_wvalid_143 && 0) begin
            write_burst_done_148 <= 1;
          end 
          if(write_burst_block_ram_wvalid_143 && (write_burst_length_147 <= 1)) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
          if(write_burst_block_ram_wvalid_143 && 0) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
          if(write_burst_block_ram_wquit_144) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_17_1 = 1;
  localparam write_burst_block_fsm_17_2 = 2;
  localparam write_burst_block_fsm_17_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
      write_burst_block_length_149 <= 0;
      write_burst_block_blocksize_150 <= 0;
      write_burst_block_done_151 <= 0;
      write_burst_block_count_152 <= 0;
    end else begin
      case(write_burst_block_fsm_17)
        write_burst_block_fsm_17_init: begin
          write_burst_block_length_149 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_150 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_151 <= 0;
          write_burst_block_count_152 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_1;
          end 
        end
        write_burst_block_fsm_17_1: begin
          if(maxi_rvalid) begin
            write_burst_block_length_149 <= write_burst_block_length_149 - 1;
            write_burst_block_done_151 <= 0;
            write_burst_block_count_152 <= write_burst_block_count_152 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_149 <= 1)) begin
            write_burst_block_done_151 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_151 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_152 == write_burst_block_blocksize_150 - 1)) begin
            write_burst_block_count_152 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_152 == write_burst_block_blocksize_150 - 1)) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_2;
          end 
          if(maxi_rvalid && (write_burst_block_length_149 <= 1)) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
          if(0) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
        end
        write_burst_block_fsm_17_2: begin
          if(maxi_rvalid) begin
            write_burst_block_length_149 <= write_burst_block_length_149 - 1;
            write_burst_block_done_151 <= 0;
            write_burst_block_count_152 <= write_burst_block_count_152 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_149 <= 1)) begin
            write_burst_block_done_151 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_151 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_152 == write_burst_block_blocksize_150 - 1)) begin
            write_burst_block_count_152 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_152 == write_burst_block_blocksize_150 - 1)) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_3;
          end 
          if(maxi_rvalid && (write_burst_block_length_149 <= 1)) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
          if(0) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
        end
        write_burst_block_fsm_17_3: begin
          if(maxi_rvalid) begin
            write_burst_block_length_149 <= write_burst_block_length_149 - 1;
            write_burst_block_done_151 <= 0;
            write_burst_block_count_152 <= write_burst_block_count_152 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_149 <= 1)) begin
            write_burst_block_done_151 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_151 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_152 == write_burst_block_blocksize_150 - 1)) begin
            write_burst_block_count_152 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_152 == write_burst_block_blocksize_150 - 1)) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_1;
          end 
          if(maxi_rvalid && (write_burst_block_length_149 <= 1)) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
          if(0) begin
            write_burst_block_fsm_17 <= write_burst_block_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_18_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_18 <= write_burst_fsm_18_init;
      write_burst_addr_157 <= 0;
      write_burst_stride_158 <= 0;
      write_burst_length_159 <= 0;
      write_burst_done_160 <= 0;
    end else begin
      case(write_burst_fsm_18)
        write_burst_fsm_18_init: begin
          write_burst_addr_157 <= _maxi_read_local_addr_buf;
          write_burst_stride_158 <= _maxi_read_local_stride_buf;
          write_burst_length_159 <= _maxi_read_local_size_buf;
          write_burst_done_160 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_18 <= write_burst_fsm_18_1;
          end 
        end
        write_burst_fsm_18_1: begin
          if(write_burst_block_ram_wvalid_155) begin
            write_burst_addr_157 <= write_burst_addr_157 + write_burst_stride_158;
            write_burst_length_159 <= write_burst_length_159 - 1;
            write_burst_done_160 <= 0;
          end 
          if(write_burst_block_ram_wvalid_155 && (write_burst_length_159 <= 1)) begin
            write_burst_done_160 <= 1;
          end 
          if(write_burst_block_ram_wvalid_155 && 0) begin
            write_burst_done_160 <= 1;
          end 
          if(write_burst_block_ram_wvalid_155 && (write_burst_length_159 <= 1)) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
          if(write_burst_block_ram_wvalid_155 && 0) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
          if(write_burst_block_ram_wquit_156) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_19_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_19 <= write_burst_fsm_19_init;
      write_burst_addr_163 <= 0;
      write_burst_stride_164 <= 0;
      write_burst_length_165 <= 0;
      write_burst_done_166 <= 0;
    end else begin
      case(write_burst_fsm_19)
        write_burst_fsm_19_init: begin
          write_burst_addr_163 <= _maxi_read_local_addr_buf;
          write_burst_stride_164 <= _maxi_read_local_stride_buf;
          write_burst_length_165 <= _maxi_read_local_size_buf;
          write_burst_done_166 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_19 <= write_burst_fsm_19_1;
          end 
        end
        write_burst_fsm_19_1: begin
          if(write_burst_block_ram_wvalid_161) begin
            write_burst_addr_163 <= write_burst_addr_163 + write_burst_stride_164;
            write_burst_length_165 <= write_burst_length_165 - 1;
            write_burst_done_166 <= 0;
          end 
          if(write_burst_block_ram_wvalid_161 && (write_burst_length_165 <= 1)) begin
            write_burst_done_166 <= 1;
          end 
          if(write_burst_block_ram_wvalid_161 && 0) begin
            write_burst_done_166 <= 1;
          end 
          if(write_burst_block_ram_wvalid_161 && (write_burst_length_165 <= 1)) begin
            write_burst_fsm_19 <= write_burst_fsm_19_init;
          end 
          if(write_burst_block_ram_wvalid_161 && 0) begin
            write_burst_fsm_19 <= write_burst_fsm_19_init;
          end 
          if(write_burst_block_ram_wquit_162) begin
            write_burst_fsm_19 <= write_burst_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_20_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_20 <= write_burst_fsm_20_init;
      write_burst_addr_169 <= 0;
      write_burst_stride_170 <= 0;
      write_burst_length_171 <= 0;
      write_burst_done_172 <= 0;
    end else begin
      case(write_burst_fsm_20)
        write_burst_fsm_20_init: begin
          write_burst_addr_169 <= _maxi_read_local_addr_buf;
          write_burst_stride_170 <= _maxi_read_local_stride_buf;
          write_burst_length_171 <= _maxi_read_local_size_buf;
          write_burst_done_172 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_20 <= write_burst_fsm_20_1;
          end 
        end
        write_burst_fsm_20_1: begin
          if(write_burst_block_ram_wvalid_167) begin
            write_burst_addr_169 <= write_burst_addr_169 + write_burst_stride_170;
            write_burst_length_171 <= write_burst_length_171 - 1;
            write_burst_done_172 <= 0;
          end 
          if(write_burst_block_ram_wvalid_167 && (write_burst_length_171 <= 1)) begin
            write_burst_done_172 <= 1;
          end 
          if(write_burst_block_ram_wvalid_167 && 0) begin
            write_burst_done_172 <= 1;
          end 
          if(write_burst_block_ram_wvalid_167 && (write_burst_length_171 <= 1)) begin
            write_burst_fsm_20 <= write_burst_fsm_20_init;
          end 
          if(write_burst_block_ram_wvalid_167 && 0) begin
            write_burst_fsm_20 <= write_burst_fsm_20_init;
          end 
          if(write_burst_block_ram_wquit_168) begin
            write_burst_fsm_20 <= write_burst_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_21_1 = 1;
  localparam write_burst_block_fsm_21_2 = 2;
  localparam write_burst_block_fsm_21_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
      write_burst_block_length_173 <= 0;
      write_burst_block_blocksize_174 <= 0;
      write_burst_block_done_175 <= 0;
      write_burst_block_count_176 <= 0;
    end else begin
      case(write_burst_block_fsm_21)
        write_burst_block_fsm_21_init: begin
          write_burst_block_length_173 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_174 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_175 <= 0;
          write_burst_block_count_176 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_1;
          end 
        end
        write_burst_block_fsm_21_1: begin
          if(maxi_rvalid) begin
            write_burst_block_length_173 <= write_burst_block_length_173 - 1;
            write_burst_block_done_175 <= 0;
            write_burst_block_count_176 <= write_burst_block_count_176 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_173 <= 1)) begin
            write_burst_block_done_175 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_175 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_176 == write_burst_block_blocksize_174 - 1)) begin
            write_burst_block_count_176 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_176 == write_burst_block_blocksize_174 - 1)) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_2;
          end 
          if(maxi_rvalid && (write_burst_block_length_173 <= 1)) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
          if(0) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
        end
        write_burst_block_fsm_21_2: begin
          if(maxi_rvalid) begin
            write_burst_block_length_173 <= write_burst_block_length_173 - 1;
            write_burst_block_done_175 <= 0;
            write_burst_block_count_176 <= write_burst_block_count_176 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_173 <= 1)) begin
            write_burst_block_done_175 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_175 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_176 == write_burst_block_blocksize_174 - 1)) begin
            write_burst_block_count_176 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_176 == write_burst_block_blocksize_174 - 1)) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_3;
          end 
          if(maxi_rvalid && (write_burst_block_length_173 <= 1)) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
          if(0) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
        end
        write_burst_block_fsm_21_3: begin
          if(maxi_rvalid) begin
            write_burst_block_length_173 <= write_burst_block_length_173 - 1;
            write_burst_block_done_175 <= 0;
            write_burst_block_count_176 <= write_burst_block_count_176 + 1;
          end 
          if(maxi_rvalid && (write_burst_block_length_173 <= 1)) begin
            write_burst_block_done_175 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_done_175 <= 1;
          end 
          if(maxi_rvalid && (write_burst_block_count_176 == write_burst_block_blocksize_174 - 1)) begin
            write_burst_block_count_176 <= 0;
          end 
          if(maxi_rvalid && (write_burst_block_count_176 == write_burst_block_blocksize_174 - 1)) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_1;
          end 
          if(maxi_rvalid && (write_burst_block_length_173 <= 1)) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
          if(0) begin
            write_burst_block_fsm_21 <= write_burst_block_fsm_21_init;
          end 
        end
      endcase
    end
  end

  localparam conv2d_2_comp_fsm_1 = 1;
  localparam conv2d_2_comp_fsm_2 = 2;
  localparam conv2d_2_comp_fsm_3 = 3;
  localparam conv2d_2_comp_fsm_4 = 4;
  localparam conv2d_2_comp_fsm_5 = 5;
  localparam conv2d_2_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      conv2d_2_comp_fsm <= conv2d_2_comp_fsm_init;
      conv2d_2_stream_act_local_0 <= 0;
      conv2d_2_stream_act_local_1 <= 0;
      conv2d_2_stream_act_local_2 <= 0;
      conv2d_2_stream_act_local_3 <= 0;
      conv2d_2_stream_act_local_4 <= 0;
      conv2d_2_stream_act_local_5 <= 0;
      conv2d_2_stream_act_local_6 <= 0;
      conv2d_2_stream_act_local_7 <= 0;
      conv2d_2_stream_act_local_8 <= 0;
      conv2d_2_stream_out_local_col <= 0;
      conv2d_2_stream_out_local_val <= 0;
      conv2d_2_col_count <= 0;
      conv2d_2_col_select <= 0;
      conv2d_2_filter_page_comp_offset_buf <= 0;
      conv2d_2_act_page_comp_offset_buf_0 <= 0;
      conv2d_2_act_page_comp_offset_buf_1 <= 0;
      conv2d_2_act_page_comp_offset_buf_2 <= 0;
      conv2d_2_out_page_comp_offset_buf <= 0;
      conv2d_2_row_count_buf <= 0;
      conv2d_2_row_select_buf <= 0;
      conv2d_2_och_count_buf <= 0;
      conv2d_2_next_stream_num_ops <= 0;
      conv2d_2_stream_pad_masks <= 0;
      conv2d_2_sync_comp_count <= 0;
    end else begin
      if(_stream_conv2d_2_sink_stop) begin
        conv2d_2_sync_comp_count <= conv2d_2_sync_comp_count + 1;
      end 
      if(control_conv2d_2 == 2) begin
        conv2d_2_sync_comp_count <= 0;
      end 
      case(conv2d_2_comp_fsm)
        conv2d_2_comp_fsm_init: begin
          if((control_conv2d_2 == 21) && !conv2d_2_skip_comp) begin
            conv2d_2_comp_fsm <= conv2d_2_comp_fsm_1;
          end 
        end
        conv2d_2_comp_fsm_1: begin
          conv2d_2_stream_act_local_0 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_0) begin
            conv2d_2_stream_act_local_0 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_0) begin
            conv2d_2_stream_act_local_0 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_1 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_1) begin
            conv2d_2_stream_act_local_1 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_1) begin
            conv2d_2_stream_act_local_1 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_2 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_2) begin
            conv2d_2_stream_act_local_2 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_2) begin
            conv2d_2_stream_act_local_2 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_3 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_0) begin
            conv2d_2_stream_act_local_3 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_0) begin
            conv2d_2_stream_act_local_3 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_4 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_1) begin
            conv2d_2_stream_act_local_4 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_1) begin
            conv2d_2_stream_act_local_4 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_5 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_2) begin
            conv2d_2_stream_act_local_5 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_2) begin
            conv2d_2_stream_act_local_5 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_6 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_0) begin
            conv2d_2_stream_act_local_6 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_0) begin
            conv2d_2_stream_act_local_6 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_7 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_1) begin
            conv2d_2_stream_act_local_7 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_1) begin
            conv2d_2_stream_act_local_7 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_act_local_8 <= 0;
          if(cparam_conv2d_2_stream_act_local_small_flags_2) begin
            conv2d_2_stream_act_local_8 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_2_stream_act_local_large_flags_2) begin
            conv2d_2_stream_act_local_8 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          conv2d_2_stream_out_local_col <= 0;
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_och_count == 0)) begin
            conv2d_2_stream_out_local_val <= 0;
          end 
          conv2d_2_col_count <= 0;
          conv2d_2_col_select <= cparam_conv2d_2_col_select_initval;
          conv2d_2_filter_page_comp_offset_buf <= conv2d_2_filter_page_comp_offset;
          conv2d_2_act_page_comp_offset_buf_0 <= conv2d_2_act_page_comp_offset_0;
          conv2d_2_act_page_comp_offset_buf_1 <= conv2d_2_act_page_comp_offset_1;
          conv2d_2_act_page_comp_offset_buf_2 <= conv2d_2_act_page_comp_offset_2;
          conv2d_2_out_page_comp_offset_buf <= conv2d_2_out_page_comp_offset;
          conv2d_2_row_count_buf <= conv2d_2_row_count;
          conv2d_2_row_select_buf <= conv2d_2_row_select;
          conv2d_2_och_count_buf <= conv2d_2_och_count;
          conv2d_2_next_stream_num_ops <= (conv2d_2_och_count >= cparam_conv2d_2_max_och_count)? cparam_conv2d_2_stream_num_ops_res : cparam_conv2d_2_stream_num_ops;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_2;
        end
        conv2d_2_comp_fsm_2: begin
          conv2d_2_stream_pad_masks <= { conv2d_2_stream_pad_mask_2_2, conv2d_2_stream_pad_mask_2_1, conv2d_2_stream_pad_mask_2_0, conv2d_2_stream_pad_mask_1_2, conv2d_2_stream_pad_mask_1_1, conv2d_2_stream_pad_mask_1_0, conv2d_2_stream_pad_mask_0_2, conv2d_2_stream_pad_mask_0_1, conv2d_2_stream_pad_mask_0_0 };
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_3;
        end
        conv2d_2_comp_fsm_3: begin
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          if(_stream_conv2d_2_stream_oready) begin
            conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
          end 
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_4;
        end
        conv2d_2_comp_fsm_4: begin
          if(!_stream_conv2d_2_source_busy) begin
            conv2d_2_comp_fsm <= conv2d_2_comp_fsm_5;
          end 
        end
        conv2d_2_comp_fsm_5: begin
          if(_stream_conv2d_2_busy) begin
            conv2d_2_comp_fsm <= conv2d_2_comp_fsm_6;
          end 
        end
        conv2d_2_comp_fsm_6: begin
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_0 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_1 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_2 : 0)) begin
            conv2d_2_stream_act_local_0 <= conv2d_2_stream_act_local_0 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_0 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_1 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_2 : 0) begin
            conv2d_2_stream_act_local_0 <= conv2d_2_stream_act_local_0 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_0 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_0) begin
            conv2d_2_stream_act_local_0 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_0) begin
            conv2d_2_stream_act_local_0 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_3 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_4 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_5 : 0)) begin
            conv2d_2_stream_act_local_1 <= conv2d_2_stream_act_local_1 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_3 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_4 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_5 : 0) begin
            conv2d_2_stream_act_local_1 <= conv2d_2_stream_act_local_1 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_1 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_1) begin
            conv2d_2_stream_act_local_1 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_1) begin
            conv2d_2_stream_act_local_1 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_6 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_7 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_8 : 0)) begin
            conv2d_2_stream_act_local_2 <= conv2d_2_stream_act_local_2 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_6 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_7 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_8 : 0) begin
            conv2d_2_stream_act_local_2 <= conv2d_2_stream_act_local_2 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_2 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_2) begin
            conv2d_2_stream_act_local_2 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_2) begin
            conv2d_2_stream_act_local_2 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_9 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_10 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_11 : 0)) begin
            conv2d_2_stream_act_local_3 <= conv2d_2_stream_act_local_3 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_9 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_10 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_11 : 0) begin
            conv2d_2_stream_act_local_3 <= conv2d_2_stream_act_local_3 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_3 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_0) begin
            conv2d_2_stream_act_local_3 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_0) begin
            conv2d_2_stream_act_local_3 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_12 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_13 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_14 : 0)) begin
            conv2d_2_stream_act_local_4 <= conv2d_2_stream_act_local_4 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_12 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_13 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_14 : 0) begin
            conv2d_2_stream_act_local_4 <= conv2d_2_stream_act_local_4 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_4 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_1) begin
            conv2d_2_stream_act_local_4 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_1) begin
            conv2d_2_stream_act_local_4 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_15 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_16 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_17 : 0)) begin
            conv2d_2_stream_act_local_5 <= conv2d_2_stream_act_local_5 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_15 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_16 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_17 : 0) begin
            conv2d_2_stream_act_local_5 <= conv2d_2_stream_act_local_5 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_5 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_2) begin
            conv2d_2_stream_act_local_5 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_2) begin
            conv2d_2_stream_act_local_5 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_18 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_19 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_20 : 0)) begin
            conv2d_2_stream_act_local_6 <= conv2d_2_stream_act_local_6 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_18 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_19 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_20 : 0) begin
            conv2d_2_stream_act_local_6 <= conv2d_2_stream_act_local_6 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_6 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_0) begin
            conv2d_2_stream_act_local_6 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_0) begin
            conv2d_2_stream_act_local_6 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_21 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_22 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_23 : 0)) begin
            conv2d_2_stream_act_local_7 <= conv2d_2_stream_act_local_7 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_21 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_22 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_23 : 0) begin
            conv2d_2_stream_act_local_7 <= conv2d_2_stream_act_local_7 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_7 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_1) begin
            conv2d_2_stream_act_local_7 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_1) begin
            conv2d_2_stream_act_local_7 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(!((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_24 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_25 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_26 : 0)) begin
            conv2d_2_stream_act_local_8 <= conv2d_2_stream_act_local_8 + cparam_conv2d_2_inc_act_laddr_small;
          end 
          if((conv2d_2_col_select == 0)? cparam_conv2d_2_inc_act_laddr_conds_24 : 
          (conv2d_2_col_select == 1)? cparam_conv2d_2_inc_act_laddr_conds_25 : 
          (conv2d_2_col_select == 2)? cparam_conv2d_2_inc_act_laddr_conds_26 : 0) begin
            conv2d_2_stream_act_local_8 <= conv2d_2_stream_act_local_8 + cparam_conv2d_2_inc_act_laddr_large;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_stream_act_local_8 <= 0;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_small_flags_2) begin
            conv2d_2_stream_act_local_8 <= cparam_conv2d_2_stream_act_local_small_offset;
          end 
          if((conv2d_2_col_count >= cparam_conv2d_2_max_col_count) && cparam_conv2d_2_stream_act_local_large_flags_2) begin
            conv2d_2_stream_act_local_8 <= cparam_conv2d_2_stream_act_local_large_offset;
          end 
          if(cparam_conv2d_2_data_stationary == 0) begin
            conv2d_2_stream_out_local_col <= conv2d_2_stream_out_local_col + conv2d_2_next_stream_num_ops;
          end 
          if((cparam_conv2d_2_data_stationary == 0) && (conv2d_2_col_count >= cparam_conv2d_2_max_col_count)) begin
            conv2d_2_stream_out_local_col <= 0;
          end 
          if(cparam_conv2d_2_data_stationary == 1) begin
            conv2d_2_stream_out_local_col <= conv2d_2_stream_out_local_col + cparam_conv2d_2_inc_out_laddr_col;
          end 
          if((cparam_conv2d_2_data_stationary == 1) && (conv2d_2_col_count >= cparam_conv2d_2_max_col_count)) begin
            conv2d_2_stream_out_local_val <= conv2d_2_stream_out_local_val + conv2d_2_next_stream_num_ops;
            conv2d_2_stream_out_local_col <= 0;
          end 
          conv2d_2_col_count <= conv2d_2_col_count + cparam_conv2d_2_stride_col_par_col;
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_col_count <= 0;
          end 
          conv2d_2_col_select <= conv2d_2_col_select + cparam_conv2d_2_stride_col_mod_filter_num;
          if(conv2d_2_col_select + cparam_conv2d_2_stride_col_mod_filter_num >= 3) begin
            conv2d_2_col_select <= conv2d_2_col_select - cparam_conv2d_2_filter_num_col_minus_stride_col_mod;
          end 
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_col_select <= cparam_conv2d_2_col_select_initval;
          end 
          conv2d_2_comp_fsm <= conv2d_2_comp_fsm_2;
          if(conv2d_2_col_count >= cparam_conv2d_2_max_col_count) begin
            conv2d_2_comp_fsm <= conv2d_2_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_20_source_pat_fsm_0_1 = 1;
  localparam _stream_conv2d_2_source_20_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_20_source_pat_fsm_0 <= _stream_conv2d_2_source_20_source_pat_fsm_0_init;
    end else begin
      case(_stream_conv2d_2_source_20_source_pat_fsm_0)
        _stream_conv2d_2_source_20_source_pat_fsm_0_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_20_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_20_source_pat_fsm_0 <= _stream_conv2d_2_source_20_source_pat_fsm_0_1;
          end 
        end
        _stream_conv2d_2_source_20_source_pat_fsm_0_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_20_source_pat_fsm_0 <= _stream_conv2d_2_source_20_source_pat_fsm_0_init;
          end 
          if((_source_stream_conv2d_2_source_20_pat_count_0 == 0) && (_source_stream_conv2d_2_source_20_pat_count_1 == 0) && (_source_stream_conv2d_2_source_20_pat_count_2 == 0) && (_source_stream_conv2d_2_source_20_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_20_source_pat_fsm_0 <= _stream_conv2d_2_source_20_source_pat_fsm_0_2;
          end 
        end
        _stream_conv2d_2_source_20_source_pat_fsm_0_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_20_source_pat_fsm_0 <= _stream_conv2d_2_source_20_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_21_source_pat_fsm_1_1 = 1;
  localparam _stream_conv2d_2_source_21_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_21_source_pat_fsm_1 <= _stream_conv2d_2_source_21_source_pat_fsm_1_init;
    end else begin
      case(_stream_conv2d_2_source_21_source_pat_fsm_1)
        _stream_conv2d_2_source_21_source_pat_fsm_1_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_21_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_21_source_pat_fsm_1 <= _stream_conv2d_2_source_21_source_pat_fsm_1_1;
          end 
        end
        _stream_conv2d_2_source_21_source_pat_fsm_1_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_21_source_pat_fsm_1 <= _stream_conv2d_2_source_21_source_pat_fsm_1_init;
          end 
          if((_source_stream_conv2d_2_source_21_pat_count_0 == 0) && (_source_stream_conv2d_2_source_21_pat_count_1 == 0) && (_source_stream_conv2d_2_source_21_pat_count_2 == 0) && (_source_stream_conv2d_2_source_21_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_21_source_pat_fsm_1 <= _stream_conv2d_2_source_21_source_pat_fsm_1_2;
          end 
        end
        _stream_conv2d_2_source_21_source_pat_fsm_1_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_21_source_pat_fsm_1 <= _stream_conv2d_2_source_21_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_22_source_pat_fsm_2_1 = 1;
  localparam _stream_conv2d_2_source_22_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_22_source_pat_fsm_2 <= _stream_conv2d_2_source_22_source_pat_fsm_2_init;
    end else begin
      case(_stream_conv2d_2_source_22_source_pat_fsm_2)
        _stream_conv2d_2_source_22_source_pat_fsm_2_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_22_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_22_source_pat_fsm_2 <= _stream_conv2d_2_source_22_source_pat_fsm_2_1;
          end 
        end
        _stream_conv2d_2_source_22_source_pat_fsm_2_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_22_source_pat_fsm_2 <= _stream_conv2d_2_source_22_source_pat_fsm_2_init;
          end 
          if((_source_stream_conv2d_2_source_22_pat_count_0 == 0) && (_source_stream_conv2d_2_source_22_pat_count_1 == 0) && (_source_stream_conv2d_2_source_22_pat_count_2 == 0) && (_source_stream_conv2d_2_source_22_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_22_source_pat_fsm_2 <= _stream_conv2d_2_source_22_source_pat_fsm_2_2;
          end 
        end
        _stream_conv2d_2_source_22_source_pat_fsm_2_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_22_source_pat_fsm_2 <= _stream_conv2d_2_source_22_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_23_source_pat_fsm_3_1 = 1;
  localparam _stream_conv2d_2_source_23_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_23_source_pat_fsm_3 <= _stream_conv2d_2_source_23_source_pat_fsm_3_init;
    end else begin
      case(_stream_conv2d_2_source_23_source_pat_fsm_3)
        _stream_conv2d_2_source_23_source_pat_fsm_3_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_23_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_23_source_pat_fsm_3 <= _stream_conv2d_2_source_23_source_pat_fsm_3_1;
          end 
        end
        _stream_conv2d_2_source_23_source_pat_fsm_3_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_23_source_pat_fsm_3 <= _stream_conv2d_2_source_23_source_pat_fsm_3_init;
          end 
          if((_source_stream_conv2d_2_source_23_pat_count_0 == 0) && (_source_stream_conv2d_2_source_23_pat_count_1 == 0) && (_source_stream_conv2d_2_source_23_pat_count_2 == 0) && (_source_stream_conv2d_2_source_23_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_23_source_pat_fsm_3 <= _stream_conv2d_2_source_23_source_pat_fsm_3_2;
          end 
        end
        _stream_conv2d_2_source_23_source_pat_fsm_3_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_23_source_pat_fsm_3 <= _stream_conv2d_2_source_23_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_24_source_pat_fsm_4_1 = 1;
  localparam _stream_conv2d_2_source_24_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_24_source_pat_fsm_4 <= _stream_conv2d_2_source_24_source_pat_fsm_4_init;
    end else begin
      case(_stream_conv2d_2_source_24_source_pat_fsm_4)
        _stream_conv2d_2_source_24_source_pat_fsm_4_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_24_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_24_source_pat_fsm_4 <= _stream_conv2d_2_source_24_source_pat_fsm_4_1;
          end 
        end
        _stream_conv2d_2_source_24_source_pat_fsm_4_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_24_source_pat_fsm_4 <= _stream_conv2d_2_source_24_source_pat_fsm_4_init;
          end 
          if((_source_stream_conv2d_2_source_24_pat_count_0 == 0) && (_source_stream_conv2d_2_source_24_pat_count_1 == 0) && (_source_stream_conv2d_2_source_24_pat_count_2 == 0) && (_source_stream_conv2d_2_source_24_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_24_source_pat_fsm_4 <= _stream_conv2d_2_source_24_source_pat_fsm_4_2;
          end 
        end
        _stream_conv2d_2_source_24_source_pat_fsm_4_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_24_source_pat_fsm_4 <= _stream_conv2d_2_source_24_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_25_source_pat_fsm_5_1 = 1;
  localparam _stream_conv2d_2_source_25_source_pat_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_25_source_pat_fsm_5 <= _stream_conv2d_2_source_25_source_pat_fsm_5_init;
    end else begin
      case(_stream_conv2d_2_source_25_source_pat_fsm_5)
        _stream_conv2d_2_source_25_source_pat_fsm_5_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_25_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_25_source_pat_fsm_5 <= _stream_conv2d_2_source_25_source_pat_fsm_5_1;
          end 
        end
        _stream_conv2d_2_source_25_source_pat_fsm_5_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_25_source_pat_fsm_5 <= _stream_conv2d_2_source_25_source_pat_fsm_5_init;
          end 
          if((_source_stream_conv2d_2_source_25_pat_count_0 == 0) && (_source_stream_conv2d_2_source_25_pat_count_1 == 0) && (_source_stream_conv2d_2_source_25_pat_count_2 == 0) && (_source_stream_conv2d_2_source_25_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_25_source_pat_fsm_5 <= _stream_conv2d_2_source_25_source_pat_fsm_5_2;
          end 
        end
        _stream_conv2d_2_source_25_source_pat_fsm_5_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_25_source_pat_fsm_5 <= _stream_conv2d_2_source_25_source_pat_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_26_source_pat_fsm_6_1 = 1;
  localparam _stream_conv2d_2_source_26_source_pat_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_26_source_pat_fsm_6 <= _stream_conv2d_2_source_26_source_pat_fsm_6_init;
    end else begin
      case(_stream_conv2d_2_source_26_source_pat_fsm_6)
        _stream_conv2d_2_source_26_source_pat_fsm_6_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_26_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_26_source_pat_fsm_6 <= _stream_conv2d_2_source_26_source_pat_fsm_6_1;
          end 
        end
        _stream_conv2d_2_source_26_source_pat_fsm_6_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_26_source_pat_fsm_6 <= _stream_conv2d_2_source_26_source_pat_fsm_6_init;
          end 
          if((_source_stream_conv2d_2_source_26_pat_count_0 == 0) && (_source_stream_conv2d_2_source_26_pat_count_1 == 0) && (_source_stream_conv2d_2_source_26_pat_count_2 == 0) && (_source_stream_conv2d_2_source_26_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_26_source_pat_fsm_6 <= _stream_conv2d_2_source_26_source_pat_fsm_6_2;
          end 
        end
        _stream_conv2d_2_source_26_source_pat_fsm_6_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_26_source_pat_fsm_6 <= _stream_conv2d_2_source_26_source_pat_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_27_source_pat_fsm_7_1 = 1;
  localparam _stream_conv2d_2_source_27_source_pat_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_27_source_pat_fsm_7 <= _stream_conv2d_2_source_27_source_pat_fsm_7_init;
    end else begin
      case(_stream_conv2d_2_source_27_source_pat_fsm_7)
        _stream_conv2d_2_source_27_source_pat_fsm_7_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_27_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_27_source_pat_fsm_7 <= _stream_conv2d_2_source_27_source_pat_fsm_7_1;
          end 
        end
        _stream_conv2d_2_source_27_source_pat_fsm_7_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_27_source_pat_fsm_7 <= _stream_conv2d_2_source_27_source_pat_fsm_7_init;
          end 
          if((_source_stream_conv2d_2_source_27_pat_count_0 == 0) && (_source_stream_conv2d_2_source_27_pat_count_1 == 0) && (_source_stream_conv2d_2_source_27_pat_count_2 == 0) && (_source_stream_conv2d_2_source_27_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_27_source_pat_fsm_7 <= _stream_conv2d_2_source_27_source_pat_fsm_7_2;
          end 
        end
        _stream_conv2d_2_source_27_source_pat_fsm_7_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_27_source_pat_fsm_7 <= _stream_conv2d_2_source_27_source_pat_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_28_source_pat_fsm_8_1 = 1;
  localparam _stream_conv2d_2_source_28_source_pat_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_28_source_pat_fsm_8 <= _stream_conv2d_2_source_28_source_pat_fsm_8_init;
    end else begin
      case(_stream_conv2d_2_source_28_source_pat_fsm_8)
        _stream_conv2d_2_source_28_source_pat_fsm_8_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_28_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_28_source_pat_fsm_8 <= _stream_conv2d_2_source_28_source_pat_fsm_8_1;
          end 
        end
        _stream_conv2d_2_source_28_source_pat_fsm_8_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_28_source_pat_fsm_8 <= _stream_conv2d_2_source_28_source_pat_fsm_8_init;
          end 
          if((_source_stream_conv2d_2_source_28_pat_count_0 == 0) && (_source_stream_conv2d_2_source_28_pat_count_1 == 0) && (_source_stream_conv2d_2_source_28_pat_count_2 == 0) && (_source_stream_conv2d_2_source_28_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_28_source_pat_fsm_8 <= _stream_conv2d_2_source_28_source_pat_fsm_8_2;
          end 
        end
        _stream_conv2d_2_source_28_source_pat_fsm_8_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_28_source_pat_fsm_8 <= _stream_conv2d_2_source_28_source_pat_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_29_source_pat_fsm_9_1 = 1;
  localparam _stream_conv2d_2_source_29_source_pat_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_29_source_pat_fsm_9 <= _stream_conv2d_2_source_29_source_pat_fsm_9_init;
    end else begin
      case(_stream_conv2d_2_source_29_source_pat_fsm_9)
        _stream_conv2d_2_source_29_source_pat_fsm_9_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_29_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_29_source_pat_fsm_9 <= _stream_conv2d_2_source_29_source_pat_fsm_9_1;
          end 
        end
        _stream_conv2d_2_source_29_source_pat_fsm_9_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_29_source_pat_fsm_9 <= _stream_conv2d_2_source_29_source_pat_fsm_9_init;
          end 
          if((_source_stream_conv2d_2_source_29_pat_count_0 == 0) && (_source_stream_conv2d_2_source_29_pat_count_1 == 0) && (_source_stream_conv2d_2_source_29_pat_count_2 == 0) && (_source_stream_conv2d_2_source_29_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_29_source_pat_fsm_9 <= _stream_conv2d_2_source_29_source_pat_fsm_9_2;
          end 
        end
        _stream_conv2d_2_source_29_source_pat_fsm_9_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_29_source_pat_fsm_9 <= _stream_conv2d_2_source_29_source_pat_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_30_source_pat_fsm_10_1 = 1;
  localparam _stream_conv2d_2_source_30_source_pat_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_30_source_pat_fsm_10 <= _stream_conv2d_2_source_30_source_pat_fsm_10_init;
    end else begin
      case(_stream_conv2d_2_source_30_source_pat_fsm_10)
        _stream_conv2d_2_source_30_source_pat_fsm_10_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_30_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_30_source_pat_fsm_10 <= _stream_conv2d_2_source_30_source_pat_fsm_10_1;
          end 
        end
        _stream_conv2d_2_source_30_source_pat_fsm_10_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_30_source_pat_fsm_10 <= _stream_conv2d_2_source_30_source_pat_fsm_10_init;
          end 
          if((_source_stream_conv2d_2_source_30_pat_count_0 == 0) && (_source_stream_conv2d_2_source_30_pat_count_1 == 0) && (_source_stream_conv2d_2_source_30_pat_count_2 == 0) && (_source_stream_conv2d_2_source_30_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_30_source_pat_fsm_10 <= _stream_conv2d_2_source_30_source_pat_fsm_10_2;
          end 
        end
        _stream_conv2d_2_source_30_source_pat_fsm_10_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_30_source_pat_fsm_10 <= _stream_conv2d_2_source_30_source_pat_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_31_source_pat_fsm_11_1 = 1;
  localparam _stream_conv2d_2_source_31_source_pat_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_31_source_pat_fsm_11 <= _stream_conv2d_2_source_31_source_pat_fsm_11_init;
    end else begin
      case(_stream_conv2d_2_source_31_source_pat_fsm_11)
        _stream_conv2d_2_source_31_source_pat_fsm_11_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_31_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_31_source_pat_fsm_11 <= _stream_conv2d_2_source_31_source_pat_fsm_11_1;
          end 
        end
        _stream_conv2d_2_source_31_source_pat_fsm_11_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_31_source_pat_fsm_11 <= _stream_conv2d_2_source_31_source_pat_fsm_11_init;
          end 
          if((_source_stream_conv2d_2_source_31_pat_count_0 == 0) && (_source_stream_conv2d_2_source_31_pat_count_1 == 0) && (_source_stream_conv2d_2_source_31_pat_count_2 == 0) && (_source_stream_conv2d_2_source_31_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_31_source_pat_fsm_11 <= _stream_conv2d_2_source_31_source_pat_fsm_11_2;
          end 
        end
        _stream_conv2d_2_source_31_source_pat_fsm_11_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_31_source_pat_fsm_11 <= _stream_conv2d_2_source_31_source_pat_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_32_source_pat_fsm_12_1 = 1;
  localparam _stream_conv2d_2_source_32_source_pat_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_32_source_pat_fsm_12 <= _stream_conv2d_2_source_32_source_pat_fsm_12_init;
    end else begin
      case(_stream_conv2d_2_source_32_source_pat_fsm_12)
        _stream_conv2d_2_source_32_source_pat_fsm_12_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_32_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_32_source_pat_fsm_12 <= _stream_conv2d_2_source_32_source_pat_fsm_12_1;
          end 
        end
        _stream_conv2d_2_source_32_source_pat_fsm_12_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_32_source_pat_fsm_12 <= _stream_conv2d_2_source_32_source_pat_fsm_12_init;
          end 
          if((_source_stream_conv2d_2_source_32_pat_count_0 == 0) && (_source_stream_conv2d_2_source_32_pat_count_1 == 0) && (_source_stream_conv2d_2_source_32_pat_count_2 == 0) && (_source_stream_conv2d_2_source_32_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_32_source_pat_fsm_12 <= _stream_conv2d_2_source_32_source_pat_fsm_12_2;
          end 
        end
        _stream_conv2d_2_source_32_source_pat_fsm_12_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_32_source_pat_fsm_12 <= _stream_conv2d_2_source_32_source_pat_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_33_source_pat_fsm_13_1 = 1;
  localparam _stream_conv2d_2_source_33_source_pat_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_33_source_pat_fsm_13 <= _stream_conv2d_2_source_33_source_pat_fsm_13_init;
    end else begin
      case(_stream_conv2d_2_source_33_source_pat_fsm_13)
        _stream_conv2d_2_source_33_source_pat_fsm_13_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_33_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_33_source_pat_fsm_13 <= _stream_conv2d_2_source_33_source_pat_fsm_13_1;
          end 
        end
        _stream_conv2d_2_source_33_source_pat_fsm_13_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_33_source_pat_fsm_13 <= _stream_conv2d_2_source_33_source_pat_fsm_13_init;
          end 
          if((_source_stream_conv2d_2_source_33_pat_count_0 == 0) && (_source_stream_conv2d_2_source_33_pat_count_1 == 0) && (_source_stream_conv2d_2_source_33_pat_count_2 == 0) && (_source_stream_conv2d_2_source_33_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_33_source_pat_fsm_13 <= _stream_conv2d_2_source_33_source_pat_fsm_13_2;
          end 
        end
        _stream_conv2d_2_source_33_source_pat_fsm_13_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_33_source_pat_fsm_13 <= _stream_conv2d_2_source_33_source_pat_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_34_source_pat_fsm_14_1 = 1;
  localparam _stream_conv2d_2_source_34_source_pat_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_34_source_pat_fsm_14 <= _stream_conv2d_2_source_34_source_pat_fsm_14_init;
    end else begin
      case(_stream_conv2d_2_source_34_source_pat_fsm_14)
        _stream_conv2d_2_source_34_source_pat_fsm_14_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_34_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_34_source_pat_fsm_14 <= _stream_conv2d_2_source_34_source_pat_fsm_14_1;
          end 
        end
        _stream_conv2d_2_source_34_source_pat_fsm_14_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_34_source_pat_fsm_14 <= _stream_conv2d_2_source_34_source_pat_fsm_14_init;
          end 
          if((_source_stream_conv2d_2_source_34_pat_count_0 == 0) && (_source_stream_conv2d_2_source_34_pat_count_1 == 0) && (_source_stream_conv2d_2_source_34_pat_count_2 == 0) && (_source_stream_conv2d_2_source_34_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_34_source_pat_fsm_14 <= _stream_conv2d_2_source_34_source_pat_fsm_14_2;
          end 
        end
        _stream_conv2d_2_source_34_source_pat_fsm_14_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_34_source_pat_fsm_14 <= _stream_conv2d_2_source_34_source_pat_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_35_source_pat_fsm_15_1 = 1;
  localparam _stream_conv2d_2_source_35_source_pat_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_35_source_pat_fsm_15 <= _stream_conv2d_2_source_35_source_pat_fsm_15_init;
    end else begin
      case(_stream_conv2d_2_source_35_source_pat_fsm_15)
        _stream_conv2d_2_source_35_source_pat_fsm_15_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_35_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_35_source_pat_fsm_15 <= _stream_conv2d_2_source_35_source_pat_fsm_15_1;
          end 
        end
        _stream_conv2d_2_source_35_source_pat_fsm_15_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_35_source_pat_fsm_15 <= _stream_conv2d_2_source_35_source_pat_fsm_15_init;
          end 
          if((_source_stream_conv2d_2_source_35_pat_count_0 == 0) && (_source_stream_conv2d_2_source_35_pat_count_1 == 0) && (_source_stream_conv2d_2_source_35_pat_count_2 == 0) && (_source_stream_conv2d_2_source_35_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_35_source_pat_fsm_15 <= _stream_conv2d_2_source_35_source_pat_fsm_15_2;
          end 
        end
        _stream_conv2d_2_source_35_source_pat_fsm_15_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_35_source_pat_fsm_15 <= _stream_conv2d_2_source_35_source_pat_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_36_source_pat_fsm_16_1 = 1;
  localparam _stream_conv2d_2_source_36_source_pat_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_36_source_pat_fsm_16 <= _stream_conv2d_2_source_36_source_pat_fsm_16_init;
    end else begin
      case(_stream_conv2d_2_source_36_source_pat_fsm_16)
        _stream_conv2d_2_source_36_source_pat_fsm_16_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_36_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_36_source_pat_fsm_16 <= _stream_conv2d_2_source_36_source_pat_fsm_16_1;
          end 
        end
        _stream_conv2d_2_source_36_source_pat_fsm_16_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_36_source_pat_fsm_16 <= _stream_conv2d_2_source_36_source_pat_fsm_16_init;
          end 
          if((_source_stream_conv2d_2_source_36_pat_count_0 == 0) && (_source_stream_conv2d_2_source_36_pat_count_1 == 0) && (_source_stream_conv2d_2_source_36_pat_count_2 == 0) && (_source_stream_conv2d_2_source_36_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_36_source_pat_fsm_16 <= _stream_conv2d_2_source_36_source_pat_fsm_16_2;
          end 
        end
        _stream_conv2d_2_source_36_source_pat_fsm_16_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_36_source_pat_fsm_16 <= _stream_conv2d_2_source_36_source_pat_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_source_37_source_pat_fsm_17_1 = 1;
  localparam _stream_conv2d_2_source_37_source_pat_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_source_37_source_pat_fsm_17 <= _stream_conv2d_2_source_37_source_pat_fsm_17_init;
    end else begin
      case(_stream_conv2d_2_source_37_source_pat_fsm_17)
        _stream_conv2d_2_source_37_source_pat_fsm_17_init: begin
          if(_stream_conv2d_2_source_start && _stream_conv2d_2_source_37_source_mode & 5'b10 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_37_source_pat_fsm_17 <= _stream_conv2d_2_source_37_source_pat_fsm_17_1;
          end 
        end
        _stream_conv2d_2_source_37_source_pat_fsm_17_1: begin
          if(_stream_conv2d_2_source_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_37_source_pat_fsm_17 <= _stream_conv2d_2_source_37_source_pat_fsm_17_init;
          end 
          if((_source_stream_conv2d_2_source_37_pat_count_0 == 0) && (_source_stream_conv2d_2_source_37_pat_count_1 == 0) && (_source_stream_conv2d_2_source_37_pat_count_2 == 0) && (_source_stream_conv2d_2_source_37_pat_count_3 == 0) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_37_source_pat_fsm_17 <= _stream_conv2d_2_source_37_source_pat_fsm_17_2;
          end 
        end
        _stream_conv2d_2_source_37_source_pat_fsm_17_2: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_source_37_source_pat_fsm_17 <= _stream_conv2d_2_source_37_source_pat_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_2_sink_50_sink_fsm_18_1 = 1;
  localparam _stream_conv2d_2_sink_50_sink_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_2_sink_50_sink_fsm_18 <= _stream_conv2d_2_sink_50_sink_fsm_18_init;
    end else begin
      case(_stream_conv2d_2_sink_50_sink_fsm_18)
        _stream_conv2d_2_sink_50_sink_fsm_18_init: begin
          if(_stream_conv2d_2_sink_start && _stream_conv2d_2_sink_50_sink_mode & 5'b1 && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_sink_50_sink_fsm_18 <= _stream_conv2d_2_sink_50_sink_fsm_18_1;
          end 
        end
        _stream_conv2d_2_sink_50_sink_fsm_18_1: begin
          if(_stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_sink_50_sink_fsm_18 <= _stream_conv2d_2_sink_50_sink_fsm_18_2;
          end 
        end
        _stream_conv2d_2_sink_50_sink_fsm_18_2: begin
          if(stream_conv2d_2_sink_51_data && (_stream_conv2d_2_sink_50_sink_count == 1) && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_sink_50_sink_fsm_18 <= _stream_conv2d_2_sink_50_sink_fsm_18_init;
          end 
          if(_stream_conv2d_2_sink_stop && _stream_conv2d_2_stream_oready) begin
            _stream_conv2d_2_sink_50_sink_fsm_18 <= _stream_conv2d_2_sink_50_sink_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
      _maxi_write_cont <= 0;
    end else begin
      case(_maxi_write_req_fsm)
        _maxi_write_req_fsm_init: begin
          if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_1;
          end 
        end
        _maxi_write_req_fsm_1: begin
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6)) begin
            _maxi_write_cont <= 1;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6) && (_maxi_write_global_size == 0)) begin
            _maxi_write_cont <= 0;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (outstanding_wcount_0 < 6)) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_data_fsm_1 = 1;
  localparam _maxi_write_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
    end else begin
      case(_maxi_write_data_fsm)
        _maxi_write_data_fsm_init: begin
          if(_maxi_write_data_idle && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(_maxi_write_data_idle && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
        end
        _maxi_write_data_fsm_1: begin
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
        end
        _maxi_write_data_fsm_2: begin
          if((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_878 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)) && read_burst_rlast_879) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_969 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0)) && read_burst_rlast_970) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_22_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_22 <= read_burst_fsm_22_init;
      read_burst_addr_875 <= 0;
      read_burst_stride_876 <= 0;
      read_burst_length_877 <= 0;
      read_burst_rvalid_878 <= 0;
      read_burst_rlast_879 <= 0;
    end else begin
      case(read_burst_fsm_22)
        read_burst_fsm_22_init: begin
          read_burst_addr_875 <= _maxi_write_local_addr_buf;
          read_burst_stride_876 <= _maxi_write_local_stride_buf;
          read_burst_length_877 <= _maxi_write_size_buf;
          read_burst_rvalid_878 <= 0;
          read_burst_rlast_879 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 1) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_22 <= read_burst_fsm_22_1;
          end 
        end
        read_burst_fsm_22_1: begin
          if((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0) && (read_burst_length_877 > 0)) begin
            read_burst_addr_875 <= read_burst_addr_875 + read_burst_stride_876;
            read_burst_length_877 <= read_burst_length_877 - 1;
            read_burst_rvalid_878 <= 1;
          end 
          if((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0) && (read_burst_length_877 <= 1)) begin
            read_burst_rlast_879 <= 1;
          end 
          if(read_burst_rlast_879 && read_burst_rvalid_878 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_878 <= 0;
            read_burst_rlast_879 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_878 <= 0;
            read_burst_rlast_879 <= 0;
          end 
          if(read_burst_rlast_879 && read_burst_rvalid_878 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_22 <= read_burst_fsm_22_init;
          end 
          if(0) begin
            read_burst_fsm_22 <= read_burst_fsm_22_init;
          end 
        end
      endcase
    end
  end

  localparam control_celu_3_1 = 1;
  localparam control_celu_3_2 = 2;
  localparam control_celu_3_3 = 3;
  localparam control_celu_3_4 = 4;
  localparam control_celu_3_5 = 5;
  localparam control_celu_3_6 = 6;
  localparam control_celu_3_7 = 7;
  localparam control_celu_3_8 = 8;
  localparam control_celu_3_9 = 9;
  localparam control_celu_3_10 = 10;
  localparam control_celu_3_11 = 11;
  localparam control_celu_3_12 = 12;
  localparam control_celu_3_13 = 13;
  localparam control_celu_3_14 = 14;
  localparam control_celu_3_15 = 15;
  localparam control_celu_3_16 = 16;
  localparam control_celu_3_17 = 17;
  localparam control_celu_3_18 = 18;
  localparam control_celu_3_19 = 19;
  localparam control_celu_3_20 = 20;
  localparam control_celu_3_21 = 21;
  localparam control_celu_3_22 = 22;
  localparam control_celu_3_23 = 23;

  always @(posedge CLK) begin
    if(RST) begin
      control_celu_3 <= control_celu_3_init;
      _control_celu_3_called <= 0;
      celu_3_out_gaddr <= 0;
      celu_3_comp_count <= 0;
      celu_3_arg_gaddr_offset_0_0 <= 0;
      celu_3_arg_gaddr_offset_0_1 <= 0;
      celu_3_arg_gaddr_offset_0_2 <= 0;
      celu_3_arg_gaddr_offset_0_3 <= 0;
      celu_3_arg_trip_count_0_0 <= 0;
      celu_3_arg_trip_count_0_1 <= 0;
      celu_3_arg_trip_count_0_2 <= 0;
      celu_3_arg_trip_count_0_3 <= 0;
      celu_3_arg_repeat_count_0_0 <= 0;
      celu_3_arg_repeat_count_0_1 <= 0;
      celu_3_arg_repeat_count_0_2 <= 0;
      celu_3_arg_repeat_count_0_3 <= 0;
      celu_3_out_page <= 0;
      celu_3_out_page_comp_offset <= 0;
      celu_3_out_page_dma_offset <= 0;
      celu_3_arg_page_0 <= 0;
      celu_3_arg_page_comp_offset_0 <= 0;
      celu_3_arg_page_dma_offset_0 <= 0;
      celu_3_skip_read <= 0;
      celu_3_skip_comp <= 0;
      celu_3_skip_write <= 0;
    end else begin
      case(control_celu_3)
        control_celu_3_init: begin
          if(main_fsm == 14) begin
            _control_celu_3_called <= 1;
          end 
          if(main_fsm == 14) begin
            control_celu_3 <= control_celu_3_1;
          end 
        end
        control_celu_3_1: begin
          control_celu_3 <= control_celu_3_2;
        end
        control_celu_3_2: begin
          celu_3_out_gaddr <= 0;
          celu_3_comp_count <= 0;
          celu_3_arg_gaddr_offset_0_0 <= 0;
          celu_3_arg_gaddr_offset_0_1 <= 0;
          celu_3_arg_gaddr_offset_0_2 <= 0;
          celu_3_arg_gaddr_offset_0_3 <= 0;
          celu_3_arg_trip_count_0_0 <= 0;
          celu_3_arg_trip_count_0_1 <= 0;
          celu_3_arg_trip_count_0_2 <= 0;
          celu_3_arg_trip_count_0_3 <= 0;
          celu_3_arg_repeat_count_0_0 <= 0;
          celu_3_arg_repeat_count_0_1 <= 0;
          celu_3_arg_repeat_count_0_2 <= 0;
          celu_3_arg_repeat_count_0_3 <= 0;
          celu_3_out_page <= 0;
          celu_3_out_page_comp_offset <= 0;
          celu_3_out_page_dma_offset <= 64;
          celu_3_arg_page_0 <= 0;
          celu_3_arg_page_comp_offset_0 <= 0;
          celu_3_arg_page_dma_offset_0 <= 0;
          celu_3_skip_read <= 0;
          celu_3_skip_comp <= 0;
          celu_3_skip_write <= 1;
          control_celu_3 <= control_celu_3_3;
        end
        control_celu_3_3: begin
          control_celu_3 <= control_celu_3_4;
          if(celu_3_skip_read) begin
            control_celu_3 <= control_celu_3_12;
          end 
        end
        control_celu_3_4: begin
          control_celu_3 <= control_celu_3_5;
          if(cparam_celu_3_arg_omit_dmas_0 && !celu_3_skip_write) begin
            control_celu_3 <= control_celu_3_12;
          end 
          if(cparam_celu_3_arg_omit_dmas_0 && cparam_celu_3_arg_stride_zeros_0 && celu_3_skip_write) begin
            control_celu_3 <= control_celu_3_8;
          end 
        end
        control_celu_3_5: begin
          if(_maxi_read_req_idle) begin
            control_celu_3 <= control_celu_3_6;
          end 
        end
        control_celu_3_6: begin
          if(_maxi_read_idle) begin
            control_celu_3 <= control_celu_3_7;
          end 
        end
        control_celu_3_7: begin
          control_celu_3 <= control_celu_3_8;
        end
        control_celu_3_8: begin
          control_celu_3 <= control_celu_3_9;
          if(!cparam_celu_3_arg_stride_zeros_0) begin
            control_celu_3 <= control_celu_3_12;
          end 
        end
        control_celu_3_9: begin
          if(_maxi_read_req_idle) begin
            control_celu_3 <= control_celu_3_10;
          end 
        end
        control_celu_3_10: begin
          if(_maxi_read_idle) begin
            control_celu_3 <= control_celu_3_11;
          end 
        end
        control_celu_3_11: begin
          control_celu_3 <= control_celu_3_12;
        end
        control_celu_3_12: begin
          if(!_stream_celu_3_source_busy) begin
            control_celu_3 <= control_celu_3_13;
          end 
          if(celu_3_skip_comp) begin
            control_celu_3 <= control_celu_3_17;
          end 
        end
        control_celu_3_13: begin
          control_celu_3 <= control_celu_3_14;
          control_celu_3 <= control_celu_3_14;
          if(_stream_celu_3_stream_oready) begin
            control_celu_3 <= control_celu_3_14;
          end 
          control_celu_3 <= control_celu_3_14;
        end
        control_celu_3_14: begin
          if(_maxi_write_idle) begin
            control_celu_3 <= control_celu_3_15;
          end 
        end
        control_celu_3_15: begin
          control_celu_3 <= control_celu_3_16;
        end
        control_celu_3_16: begin
          if(_stream_celu_3_busy) begin
            control_celu_3 <= control_celu_3_17;
          end 
        end
        control_celu_3_17: begin
          if(!_stream_celu_3_busy) begin
            control_celu_3 <= control_celu_3_18;
          end 
          if(!celu_3_skip_comp) begin
            control_celu_3 <= control_celu_3_18;
          end 
        end
        control_celu_3_18: begin
          control_celu_3 <= control_celu_3_19;
          if(celu_3_skip_write) begin
            control_celu_3 <= control_celu_3_21;
          end 
        end
        control_celu_3_19: begin
          if(_maxi_write_req_idle) begin
            control_celu_3 <= control_celu_3_20;
          end 
        end
        control_celu_3_20: begin
          control_celu_3 <= control_celu_3_21;
        end
        control_celu_3_21: begin
          celu_3_comp_count <= celu_3_comp_count + 1;
          if(!celu_3_skip_write) begin
            celu_3_out_gaddr <= celu_3_out_gaddr + cparam_celu_3_addr_inc;
          end 
          celu_3_arg_repeat_count_0_2 <= celu_3_arg_repeat_count_0_2 + 1;
          if(celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) begin
            celu_3_arg_repeat_count_0_2 <= 0;
            celu_3_arg_trip_count_0_2 <= celu_3_arg_trip_count_0_2 + 1;
            celu_3_arg_gaddr_offset_0_2 <= celu_3_arg_gaddr_offset_0_2 + cparam_celu_3_arg_addr_incs_2;
          end 
          if((celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) && (celu_3_arg_trip_count_0_2 == cparam_celu_3_arg_trip_sizes_2 - 1)) begin
            celu_3_arg_trip_count_0_2 <= 0;
            celu_3_arg_gaddr_offset_0_2 <= 0;
          end 
          if((celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) && (celu_3_arg_trip_count_0_2 == cparam_celu_3_arg_trip_sizes_2 - 1)) begin
            celu_3_arg_repeat_count_0_1 <= celu_3_arg_repeat_count_0_1 + 1;
          end 
          if((celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) && (celu_3_arg_trip_count_0_2 == cparam_celu_3_arg_trip_sizes_2 - 1) && (celu_3_arg_repeat_count_0_1 == cparam_celu_3_arg_repeat_sizes_1 - 1)) begin
            celu_3_arg_repeat_count_0_1 <= 0;
            celu_3_arg_trip_count_0_1 <= celu_3_arg_trip_count_0_1 + 1;
            celu_3_arg_gaddr_offset_0_1 <= celu_3_arg_gaddr_offset_0_1 + cparam_celu_3_arg_addr_incs_1;
          end 
          if((celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) && (celu_3_arg_trip_count_0_2 == cparam_celu_3_arg_trip_sizes_2 - 1) && (celu_3_arg_repeat_count_0_1 == cparam_celu_3_arg_repeat_sizes_1 - 1) && (celu_3_arg_trip_count_0_1 == cparam_celu_3_arg_trip_sizes_1 - 1)) begin
            celu_3_arg_trip_count_0_1 <= 0;
            celu_3_arg_gaddr_offset_0_1 <= 0;
          end 
          if((celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) && (celu_3_arg_trip_count_0_2 == cparam_celu_3_arg_trip_sizes_2 - 1) && (celu_3_arg_repeat_count_0_1 == cparam_celu_3_arg_repeat_sizes_1 - 1) && (celu_3_arg_trip_count_0_1 == cparam_celu_3_arg_trip_sizes_1 - 1)) begin
            celu_3_arg_repeat_count_0_0 <= celu_3_arg_repeat_count_0_0 + 1;
          end 
          if((celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) && (celu_3_arg_trip_count_0_2 == cparam_celu_3_arg_trip_sizes_2 - 1) && (celu_3_arg_repeat_count_0_1 == cparam_celu_3_arg_repeat_sizes_1 - 1) && (celu_3_arg_trip_count_0_1 == cparam_celu_3_arg_trip_sizes_1 - 1) && (celu_3_arg_repeat_count_0_0 == cparam_celu_3_arg_repeat_sizes_0 - 1)) begin
            celu_3_arg_repeat_count_0_0 <= 0;
            celu_3_arg_trip_count_0_0 <= celu_3_arg_trip_count_0_0 + 1;
            celu_3_arg_gaddr_offset_0_0 <= celu_3_arg_gaddr_offset_0_0 + cparam_celu_3_arg_addr_incs_0;
          end 
          if((celu_3_arg_repeat_count_0_2 == cparam_celu_3_arg_repeat_sizes_2 - 1) && (celu_3_arg_trip_count_0_2 == cparam_celu_3_arg_trip_sizes_2 - 1) && (celu_3_arg_repeat_count_0_1 == cparam_celu_3_arg_repeat_sizes_1 - 1) && (celu_3_arg_trip_count_0_1 == cparam_celu_3_arg_trip_sizes_1 - 1) && (celu_3_arg_repeat_count_0_0 == cparam_celu_3_arg_repeat_sizes_0 - 1) && (celu_3_arg_trip_count_0_0 == cparam_celu_3_arg_trip_sizes_0 - 1)) begin
            celu_3_arg_trip_count_0_0 <= 0;
            celu_3_arg_gaddr_offset_0_0 <= 0;
          end 
          if(!celu_3_arg_page_0 && !cparam_celu_3_arg_omit_dmas_0) begin
            celu_3_arg_page_comp_offset_0 <= 64;
            celu_3_arg_page_dma_offset_0 <= 64;
            celu_3_arg_page_0 <= 1;
          end 
          if(celu_3_arg_page_0 && !cparam_celu_3_arg_omit_dmas_0) begin
            celu_3_arg_page_comp_offset_0 <= 0;
            celu_3_arg_page_dma_offset_0 <= 0;
            celu_3_arg_page_0 <= 0;
          end 
          if(!celu_3_out_page) begin
            celu_3_out_page_comp_offset <= 64;
            celu_3_out_page_dma_offset <= 0;
            celu_3_out_page <= 1;
          end 
          if(celu_3_out_page) begin
            celu_3_out_page_comp_offset <= 0;
            celu_3_out_page_dma_offset <= 64;
            celu_3_out_page <= 0;
          end 
          celu_3_skip_write <= 0;
          if(celu_3_comp_count == cparam_celu_3_num_comp - 1) begin
            celu_3_skip_read <= 1;
            celu_3_skip_comp <= 1;
          end 
          if(celu_3_comp_count < cparam_celu_3_num_comp) begin
            control_celu_3 <= control_celu_3_3;
          end 
          if(celu_3_comp_count == cparam_celu_3_num_comp) begin
            control_celu_3 <= control_celu_3_22;
          end 
        end
        control_celu_3_22: begin
          if(_maxi_write_idle && (outstanding_wcount_0 == 0)) begin
            control_celu_3 <= control_celu_3_23;
          end 
        end
        control_celu_3_23: begin
          if(main_fsm == 17) begin
            _control_celu_3_called <= 0;
          end 
          if(main_fsm == 17) begin
            control_celu_3 <= control_celu_3_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_23_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_23 <= write_burst_fsm_23_init;
      write_burst_addr_885 <= 0;
      write_burst_stride_886 <= 0;
      write_burst_length_887 <= 0;
      write_burst_done_888 <= 0;
    end else begin
      case(write_burst_fsm_23)
        write_burst_fsm_23_init: begin
          write_burst_addr_885 <= _maxi_read_local_addr_buf;
          write_burst_stride_886 <= _maxi_read_local_stride_buf;
          write_burst_length_887 <= _maxi_read_local_size_buf;
          write_burst_done_888 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_23 <= write_burst_fsm_23_1;
          end 
        end
        write_burst_fsm_23_1: begin
          if(maxi_rvalid) begin
            write_burst_addr_885 <= write_burst_addr_885 + write_burst_stride_886;
            write_burst_length_887 <= write_burst_length_887 - 1;
            write_burst_done_888 <= 0;
          end 
          if(maxi_rvalid && (write_burst_length_887 <= 1)) begin
            write_burst_done_888 <= 1;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_done_888 <= 1;
          end 
          if(maxi_rvalid && (write_burst_length_887 <= 1)) begin
            write_burst_fsm_23 <= write_burst_fsm_23_init;
          end 
          if(maxi_rvalid && 0) begin
            write_burst_fsm_23 <= write_burst_fsm_23_init;
          end 
          if(0) begin
            write_burst_fsm_23 <= write_burst_fsm_23_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_celu_3_source_1_source_fsm_0_1 = 1;
  localparam _stream_celu_3_source_1_source_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_celu_3_source_1_source_fsm_0 <= _stream_celu_3_source_1_source_fsm_0_init;
    end else begin
      case(_stream_celu_3_source_1_source_fsm_0)
        _stream_celu_3_source_1_source_fsm_0_init: begin
          if(_stream_celu_3_source_start && _stream_celu_3_source_1_source_mode & 5'b1 && _stream_celu_3_stream_oready) begin
            _stream_celu_3_source_1_source_fsm_0 <= _stream_celu_3_source_1_source_fsm_0_1;
          end 
        end
        _stream_celu_3_source_1_source_fsm_0_1: begin
          if(_stream_celu_3_stream_oready) begin
            _stream_celu_3_source_1_source_fsm_0 <= _stream_celu_3_source_1_source_fsm_0_2;
          end 
        end
        _stream_celu_3_source_1_source_fsm_0_2: begin
          if((_stream_celu_3_source_1_source_count == 1) && _stream_celu_3_stream_oready) begin
            _stream_celu_3_source_1_source_fsm_0 <= _stream_celu_3_source_1_source_fsm_0_init;
          end 
          if(_stream_celu_3_source_stop && _stream_celu_3_stream_oready) begin
            _stream_celu_3_source_1_source_fsm_0 <= _stream_celu_3_source_1_source_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_celu_3_sink_2_sink_fsm_1_1 = 1;
  localparam _stream_celu_3_sink_2_sink_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_celu_3_sink_2_sink_fsm_1 <= _stream_celu_3_sink_2_sink_fsm_1_init;
    end else begin
      case(_stream_celu_3_sink_2_sink_fsm_1)
        _stream_celu_3_sink_2_sink_fsm_1_init: begin
          if(_stream_celu_3_sink_start && _stream_celu_3_sink_2_sink_mode & 5'b1 && _stream_celu_3_stream_oready) begin
            _stream_celu_3_sink_2_sink_fsm_1 <= _stream_celu_3_sink_2_sink_fsm_1_1;
          end 
        end
        _stream_celu_3_sink_2_sink_fsm_1_1: begin
          if(_stream_celu_3_stream_oready) begin
            _stream_celu_3_sink_2_sink_fsm_1 <= _stream_celu_3_sink_2_sink_fsm_1_2;
          end 
        end
        _stream_celu_3_sink_2_sink_fsm_1_2: begin
          if((_stream_celu_3_sink_2_sink_count == 1) && _stream_celu_3_stream_oready) begin
            _stream_celu_3_sink_2_sink_fsm_1 <= _stream_celu_3_sink_2_sink_fsm_1_init;
          end 
          if(_stream_celu_3_sink_stop && _stream_celu_3_stream_oready) begin
            _stream_celu_3_sink_2_sink_fsm_1 <= _stream_celu_3_sink_2_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_24_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_24 <= read_burst_fsm_24_init;
      read_burst_addr_966 <= 0;
      read_burst_stride_967 <= 0;
      read_burst_length_968 <= 0;
      read_burst_rvalid_969 <= 0;
      read_burst_rlast_970 <= 0;
    end else begin
      case(read_burst_fsm_24)
        read_burst_fsm_24_init: begin
          read_burst_addr_966 <= _maxi_write_local_addr_buf;
          read_burst_stride_967 <= _maxi_write_local_stride_buf;
          read_burst_length_968 <= _maxi_write_size_buf;
          read_burst_rvalid_969 <= 0;
          read_burst_rlast_970 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 2) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_24 <= read_burst_fsm_24_1;
          end 
        end
        read_burst_fsm_24_1: begin
          if((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0) && (read_burst_length_968 > 0)) begin
            read_burst_addr_966 <= read_burst_addr_966 + read_burst_stride_967;
            read_burst_length_968 <= read_burst_length_968 - 1;
            read_burst_rvalid_969 <= 1;
          end 
          if((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0) && (read_burst_length_968 <= 1)) begin
            read_burst_rlast_970 <= 1;
          end 
          if(read_burst_rlast_970 && read_burst_rvalid_969 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_969 <= 0;
            read_burst_rlast_970 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_969 <= 0;
            read_burst_rlast_970 <= 0;
          end 
          if(read_burst_rlast_970 && read_burst_rvalid_969 && ((maxi_wready || !maxi_wvalid) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_24 <= read_burst_fsm_24_init;
          end 
          if(0) begin
            read_burst_fsm_24 <= read_burst_fsm_24_init;
          end 
        end
      endcase
    end
  end


endmodule



module _maxi_read_req_fifo
(
  input CLK,
  input RST,
  input _maxi_read_req_fifo_enq,
  input [137-1:0] _maxi_read_req_fifo_wdata,
  output _maxi_read_req_fifo_full,
  output _maxi_read_req_fifo_almost_full,
  input _maxi_read_req_fifo_deq,
  output [137-1:0] _maxi_read_req_fifo_rdata,
  output _maxi_read_req_fifo_empty,
  output _maxi_read_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_read_req_fifo_full = is_full;
  assign _maxi_read_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_read_req_fifo_empty = is_empty;
  assign _maxi_read_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_read_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_read_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_read_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _maxi_write_req_fifo
(
  input CLK,
  input RST,
  input _maxi_write_req_fifo_enq,
  input [137-1:0] _maxi_write_req_fifo_wdata,
  output _maxi_write_req_fifo_full,
  output _maxi_write_req_fifo_almost_full,
  input _maxi_write_req_fifo_deq,
  output [137-1:0] _maxi_write_req_fifo_rdata,
  output _maxi_write_req_fifo_empty,
  output _maxi_write_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_write_req_fifo_full = is_full;
  assign _maxi_write_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_write_req_fifo_empty = is_empty;
  assign _maxi_write_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_write_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_write_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_write_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module ram_w32_l128_id0
(
  input CLK,
  input [7-1:0] ram_w32_l128_id0_0_addr,
  output [32-1:0] ram_w32_l128_id0_0_rdata,
  input [32-1:0] ram_w32_l128_id0_0_wdata,
  input ram_w32_l128_id0_0_wenable,
  input ram_w32_l128_id0_0_enable,
  input [7-1:0] ram_w32_l128_id0_1_addr,
  output [32-1:0] ram_w32_l128_id0_1_rdata,
  input [32-1:0] ram_w32_l128_id0_1_wdata,
  input ram_w32_l128_id0_1_wenable,
  input ram_w32_l128_id0_1_enable
);

  reg [32-1:0] ram_w32_l128_id0_0_rdata_out;
  assign ram_w32_l128_id0_0_rdata = ram_w32_l128_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id0_1_rdata_out;
  assign ram_w32_l128_id0_1_rdata = ram_w32_l128_id0_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id0_0_enable) begin
      if(ram_w32_l128_id0_0_wenable) begin
        mem[ram_w32_l128_id0_0_addr] <= ram_w32_l128_id0_0_wdata;
        ram_w32_l128_id0_0_rdata_out <= ram_w32_l128_id0_0_wdata;
      end else begin
        ram_w32_l128_id0_0_rdata_out <= mem[ram_w32_l128_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id0_1_enable) begin
      if(ram_w32_l128_id0_1_wenable) begin
        mem[ram_w32_l128_id0_1_addr] <= ram_w32_l128_id0_1_wdata;
        ram_w32_l128_id0_1_rdata_out <= ram_w32_l128_id0_1_wdata;
      end else begin
        ram_w32_l128_id0_1_rdata_out <= mem[ram_w32_l128_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id1
(
  input CLK,
  input [7-1:0] ram_w32_l128_id1_0_addr,
  output [32-1:0] ram_w32_l128_id1_0_rdata,
  input [32-1:0] ram_w32_l128_id1_0_wdata,
  input ram_w32_l128_id1_0_wenable,
  input ram_w32_l128_id1_0_enable,
  input [7-1:0] ram_w32_l128_id1_1_addr,
  output [32-1:0] ram_w32_l128_id1_1_rdata,
  input [32-1:0] ram_w32_l128_id1_1_wdata,
  input ram_w32_l128_id1_1_wenable,
  input ram_w32_l128_id1_1_enable
);

  reg [32-1:0] ram_w32_l128_id1_0_rdata_out;
  assign ram_w32_l128_id1_0_rdata = ram_w32_l128_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id1_1_rdata_out;
  assign ram_w32_l128_id1_1_rdata = ram_w32_l128_id1_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id1_0_enable) begin
      if(ram_w32_l128_id1_0_wenable) begin
        mem[ram_w32_l128_id1_0_addr] <= ram_w32_l128_id1_0_wdata;
        ram_w32_l128_id1_0_rdata_out <= ram_w32_l128_id1_0_wdata;
      end else begin
        ram_w32_l128_id1_0_rdata_out <= mem[ram_w32_l128_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id1_1_enable) begin
      if(ram_w32_l128_id1_1_wenable) begin
        mem[ram_w32_l128_id1_1_addr] <= ram_w32_l128_id1_1_wdata;
        ram_w32_l128_id1_1_rdata_out <= ram_w32_l128_id1_1_wdata;
      end else begin
        ram_w32_l128_id1_1_rdata_out <= mem[ram_w32_l128_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id2
(
  input CLK,
  input [7-1:0] ram_w32_l128_id2_0_addr,
  output [32-1:0] ram_w32_l128_id2_0_rdata,
  input [32-1:0] ram_w32_l128_id2_0_wdata,
  input ram_w32_l128_id2_0_wenable,
  input ram_w32_l128_id2_0_enable,
  input [7-1:0] ram_w32_l128_id2_1_addr,
  output [32-1:0] ram_w32_l128_id2_1_rdata,
  input [32-1:0] ram_w32_l128_id2_1_wdata,
  input ram_w32_l128_id2_1_wenable,
  input ram_w32_l128_id2_1_enable
);

  reg [32-1:0] ram_w32_l128_id2_0_rdata_out;
  assign ram_w32_l128_id2_0_rdata = ram_w32_l128_id2_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id2_1_rdata_out;
  assign ram_w32_l128_id2_1_rdata = ram_w32_l128_id2_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id2_0_enable) begin
      if(ram_w32_l128_id2_0_wenable) begin
        mem[ram_w32_l128_id2_0_addr] <= ram_w32_l128_id2_0_wdata;
        ram_w32_l128_id2_0_rdata_out <= ram_w32_l128_id2_0_wdata;
      end else begin
        ram_w32_l128_id2_0_rdata_out <= mem[ram_w32_l128_id2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id2_1_enable) begin
      if(ram_w32_l128_id2_1_wenable) begin
        mem[ram_w32_l128_id2_1_addr] <= ram_w32_l128_id2_1_wdata;
        ram_w32_l128_id2_1_rdata_out <= ram_w32_l128_id2_1_wdata;
      end else begin
        ram_w32_l128_id2_1_rdata_out <= mem[ram_w32_l128_id2_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id3
(
  input CLK,
  input [7-1:0] ram_w32_l128_id3_0_addr,
  output [32-1:0] ram_w32_l128_id3_0_rdata,
  input [32-1:0] ram_w32_l128_id3_0_wdata,
  input ram_w32_l128_id3_0_wenable,
  input ram_w32_l128_id3_0_enable,
  input [7-1:0] ram_w32_l128_id3_1_addr,
  output [32-1:0] ram_w32_l128_id3_1_rdata,
  input [32-1:0] ram_w32_l128_id3_1_wdata,
  input ram_w32_l128_id3_1_wenable,
  input ram_w32_l128_id3_1_enable
);

  reg [32-1:0] ram_w32_l128_id3_0_rdata_out;
  assign ram_w32_l128_id3_0_rdata = ram_w32_l128_id3_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id3_1_rdata_out;
  assign ram_w32_l128_id3_1_rdata = ram_w32_l128_id3_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id3_0_enable) begin
      if(ram_w32_l128_id3_0_wenable) begin
        mem[ram_w32_l128_id3_0_addr] <= ram_w32_l128_id3_0_wdata;
        ram_w32_l128_id3_0_rdata_out <= ram_w32_l128_id3_0_wdata;
      end else begin
        ram_w32_l128_id3_0_rdata_out <= mem[ram_w32_l128_id3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id3_1_enable) begin
      if(ram_w32_l128_id3_1_wenable) begin
        mem[ram_w32_l128_id3_1_addr] <= ram_w32_l128_id3_1_wdata;
        ram_w32_l128_id3_1_rdata_out <= ram_w32_l128_id3_1_wdata;
      end else begin
        ram_w32_l128_id3_1_rdata_out <= mem[ram_w32_l128_id3_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id4
(
  input CLK,
  input [7-1:0] ram_w32_l128_id4_0_addr,
  output [32-1:0] ram_w32_l128_id4_0_rdata,
  input [32-1:0] ram_w32_l128_id4_0_wdata,
  input ram_w32_l128_id4_0_wenable,
  input ram_w32_l128_id4_0_enable,
  input [7-1:0] ram_w32_l128_id4_1_addr,
  output [32-1:0] ram_w32_l128_id4_1_rdata,
  input [32-1:0] ram_w32_l128_id4_1_wdata,
  input ram_w32_l128_id4_1_wenable,
  input ram_w32_l128_id4_1_enable
);

  reg [32-1:0] ram_w32_l128_id4_0_rdata_out;
  assign ram_w32_l128_id4_0_rdata = ram_w32_l128_id4_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id4_1_rdata_out;
  assign ram_w32_l128_id4_1_rdata = ram_w32_l128_id4_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id4_0_enable) begin
      if(ram_w32_l128_id4_0_wenable) begin
        mem[ram_w32_l128_id4_0_addr] <= ram_w32_l128_id4_0_wdata;
        ram_w32_l128_id4_0_rdata_out <= ram_w32_l128_id4_0_wdata;
      end else begin
        ram_w32_l128_id4_0_rdata_out <= mem[ram_w32_l128_id4_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id4_1_enable) begin
      if(ram_w32_l128_id4_1_wenable) begin
        mem[ram_w32_l128_id4_1_addr] <= ram_w32_l128_id4_1_wdata;
        ram_w32_l128_id4_1_rdata_out <= ram_w32_l128_id4_1_wdata;
      end else begin
        ram_w32_l128_id4_1_rdata_out <= mem[ram_w32_l128_id4_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id5
(
  input CLK,
  input [7-1:0] ram_w32_l128_id5_0_addr,
  output [32-1:0] ram_w32_l128_id5_0_rdata,
  input [32-1:0] ram_w32_l128_id5_0_wdata,
  input ram_w32_l128_id5_0_wenable,
  input ram_w32_l128_id5_0_enable,
  input [7-1:0] ram_w32_l128_id5_1_addr,
  output [32-1:0] ram_w32_l128_id5_1_rdata,
  input [32-1:0] ram_w32_l128_id5_1_wdata,
  input ram_w32_l128_id5_1_wenable,
  input ram_w32_l128_id5_1_enable
);

  reg [32-1:0] ram_w32_l128_id5_0_rdata_out;
  assign ram_w32_l128_id5_0_rdata = ram_w32_l128_id5_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id5_1_rdata_out;
  assign ram_w32_l128_id5_1_rdata = ram_w32_l128_id5_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id5_0_enable) begin
      if(ram_w32_l128_id5_0_wenable) begin
        mem[ram_w32_l128_id5_0_addr] <= ram_w32_l128_id5_0_wdata;
        ram_w32_l128_id5_0_rdata_out <= ram_w32_l128_id5_0_wdata;
      end else begin
        ram_w32_l128_id5_0_rdata_out <= mem[ram_w32_l128_id5_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id5_1_enable) begin
      if(ram_w32_l128_id5_1_wenable) begin
        mem[ram_w32_l128_id5_1_addr] <= ram_w32_l128_id5_1_wdata;
        ram_w32_l128_id5_1_rdata_out <= ram_w32_l128_id5_1_wdata;
      end else begin
        ram_w32_l128_id5_1_rdata_out <= mem[ram_w32_l128_id5_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id6
(
  input CLK,
  input [7-1:0] ram_w32_l128_id6_0_addr,
  output [32-1:0] ram_w32_l128_id6_0_rdata,
  input [32-1:0] ram_w32_l128_id6_0_wdata,
  input ram_w32_l128_id6_0_wenable,
  input ram_w32_l128_id6_0_enable,
  input [7-1:0] ram_w32_l128_id6_1_addr,
  output [32-1:0] ram_w32_l128_id6_1_rdata,
  input [32-1:0] ram_w32_l128_id6_1_wdata,
  input ram_w32_l128_id6_1_wenable,
  input ram_w32_l128_id6_1_enable
);

  reg [32-1:0] ram_w32_l128_id6_0_rdata_out;
  assign ram_w32_l128_id6_0_rdata = ram_w32_l128_id6_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id6_1_rdata_out;
  assign ram_w32_l128_id6_1_rdata = ram_w32_l128_id6_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id6_0_enable) begin
      if(ram_w32_l128_id6_0_wenable) begin
        mem[ram_w32_l128_id6_0_addr] <= ram_w32_l128_id6_0_wdata;
        ram_w32_l128_id6_0_rdata_out <= ram_w32_l128_id6_0_wdata;
      end else begin
        ram_w32_l128_id6_0_rdata_out <= mem[ram_w32_l128_id6_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id6_1_enable) begin
      if(ram_w32_l128_id6_1_wenable) begin
        mem[ram_w32_l128_id6_1_addr] <= ram_w32_l128_id6_1_wdata;
        ram_w32_l128_id6_1_rdata_out <= ram_w32_l128_id6_1_wdata;
      end else begin
        ram_w32_l128_id6_1_rdata_out <= mem[ram_w32_l128_id6_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id7
(
  input CLK,
  input [7-1:0] ram_w32_l128_id7_0_addr,
  output [32-1:0] ram_w32_l128_id7_0_rdata,
  input [32-1:0] ram_w32_l128_id7_0_wdata,
  input ram_w32_l128_id7_0_wenable,
  input ram_w32_l128_id7_0_enable,
  input [7-1:0] ram_w32_l128_id7_1_addr,
  output [32-1:0] ram_w32_l128_id7_1_rdata,
  input [32-1:0] ram_w32_l128_id7_1_wdata,
  input ram_w32_l128_id7_1_wenable,
  input ram_w32_l128_id7_1_enable
);

  reg [32-1:0] ram_w32_l128_id7_0_rdata_out;
  assign ram_w32_l128_id7_0_rdata = ram_w32_l128_id7_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id7_1_rdata_out;
  assign ram_w32_l128_id7_1_rdata = ram_w32_l128_id7_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id7_0_enable) begin
      if(ram_w32_l128_id7_0_wenable) begin
        mem[ram_w32_l128_id7_0_addr] <= ram_w32_l128_id7_0_wdata;
        ram_w32_l128_id7_0_rdata_out <= ram_w32_l128_id7_0_wdata;
      end else begin
        ram_w32_l128_id7_0_rdata_out <= mem[ram_w32_l128_id7_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id7_1_enable) begin
      if(ram_w32_l128_id7_1_wenable) begin
        mem[ram_w32_l128_id7_1_addr] <= ram_w32_l128_id7_1_wdata;
        ram_w32_l128_id7_1_rdata_out <= ram_w32_l128_id7_1_wdata;
      end else begin
        ram_w32_l128_id7_1_rdata_out <= mem[ram_w32_l128_id7_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id8
(
  input CLK,
  input [7-1:0] ram_w32_l128_id8_0_addr,
  output [32-1:0] ram_w32_l128_id8_0_rdata,
  input [32-1:0] ram_w32_l128_id8_0_wdata,
  input ram_w32_l128_id8_0_wenable,
  input ram_w32_l128_id8_0_enable,
  input [7-1:0] ram_w32_l128_id8_1_addr,
  output [32-1:0] ram_w32_l128_id8_1_rdata,
  input [32-1:0] ram_w32_l128_id8_1_wdata,
  input ram_w32_l128_id8_1_wenable,
  input ram_w32_l128_id8_1_enable
);

  reg [32-1:0] ram_w32_l128_id8_0_rdata_out;
  assign ram_w32_l128_id8_0_rdata = ram_w32_l128_id8_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id8_1_rdata_out;
  assign ram_w32_l128_id8_1_rdata = ram_w32_l128_id8_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id8_0_enable) begin
      if(ram_w32_l128_id8_0_wenable) begin
        mem[ram_w32_l128_id8_0_addr] <= ram_w32_l128_id8_0_wdata;
        ram_w32_l128_id8_0_rdata_out <= ram_w32_l128_id8_0_wdata;
      end else begin
        ram_w32_l128_id8_0_rdata_out <= mem[ram_w32_l128_id8_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id8_1_enable) begin
      if(ram_w32_l128_id8_1_wenable) begin
        mem[ram_w32_l128_id8_1_addr] <= ram_w32_l128_id8_1_wdata;
        ram_w32_l128_id8_1_rdata_out <= ram_w32_l128_id8_1_wdata;
      end else begin
        ram_w32_l128_id8_1_rdata_out <= mem[ram_w32_l128_id8_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id9
(
  input CLK,
  input [7-1:0] ram_w32_l128_id9_0_addr,
  output [32-1:0] ram_w32_l128_id9_0_rdata,
  input [32-1:0] ram_w32_l128_id9_0_wdata,
  input ram_w32_l128_id9_0_wenable,
  input ram_w32_l128_id9_0_enable,
  input [7-1:0] ram_w32_l128_id9_1_addr,
  output [32-1:0] ram_w32_l128_id9_1_rdata,
  input [32-1:0] ram_w32_l128_id9_1_wdata,
  input ram_w32_l128_id9_1_wenable,
  input ram_w32_l128_id9_1_enable
);

  reg [32-1:0] ram_w32_l128_id9_0_rdata_out;
  assign ram_w32_l128_id9_0_rdata = ram_w32_l128_id9_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id9_1_rdata_out;
  assign ram_w32_l128_id9_1_rdata = ram_w32_l128_id9_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id9_0_enable) begin
      if(ram_w32_l128_id9_0_wenable) begin
        mem[ram_w32_l128_id9_0_addr] <= ram_w32_l128_id9_0_wdata;
        ram_w32_l128_id9_0_rdata_out <= ram_w32_l128_id9_0_wdata;
      end else begin
        ram_w32_l128_id9_0_rdata_out <= mem[ram_w32_l128_id9_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id9_1_enable) begin
      if(ram_w32_l128_id9_1_wenable) begin
        mem[ram_w32_l128_id9_1_addr] <= ram_w32_l128_id9_1_wdata;
        ram_w32_l128_id9_1_rdata_out <= ram_w32_l128_id9_1_wdata;
      end else begin
        ram_w32_l128_id9_1_rdata_out <= mem[ram_w32_l128_id9_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id10
(
  input CLK,
  input [7-1:0] ram_w32_l128_id10_0_addr,
  output [32-1:0] ram_w32_l128_id10_0_rdata,
  input [32-1:0] ram_w32_l128_id10_0_wdata,
  input ram_w32_l128_id10_0_wenable,
  input ram_w32_l128_id10_0_enable,
  input [7-1:0] ram_w32_l128_id10_1_addr,
  output [32-1:0] ram_w32_l128_id10_1_rdata,
  input [32-1:0] ram_w32_l128_id10_1_wdata,
  input ram_w32_l128_id10_1_wenable,
  input ram_w32_l128_id10_1_enable
);

  reg [32-1:0] ram_w32_l128_id10_0_rdata_out;
  assign ram_w32_l128_id10_0_rdata = ram_w32_l128_id10_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id10_1_rdata_out;
  assign ram_w32_l128_id10_1_rdata = ram_w32_l128_id10_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id10_0_enable) begin
      if(ram_w32_l128_id10_0_wenable) begin
        mem[ram_w32_l128_id10_0_addr] <= ram_w32_l128_id10_0_wdata;
        ram_w32_l128_id10_0_rdata_out <= ram_w32_l128_id10_0_wdata;
      end else begin
        ram_w32_l128_id10_0_rdata_out <= mem[ram_w32_l128_id10_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id10_1_enable) begin
      if(ram_w32_l128_id10_1_wenable) begin
        mem[ram_w32_l128_id10_1_addr] <= ram_w32_l128_id10_1_wdata;
        ram_w32_l128_id10_1_rdata_out <= ram_w32_l128_id10_1_wdata;
      end else begin
        ram_w32_l128_id10_1_rdata_out <= mem[ram_w32_l128_id10_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id11
(
  input CLK,
  input [7-1:0] ram_w32_l128_id11_0_addr,
  output [32-1:0] ram_w32_l128_id11_0_rdata,
  input [32-1:0] ram_w32_l128_id11_0_wdata,
  input ram_w32_l128_id11_0_wenable,
  input ram_w32_l128_id11_0_enable,
  input [7-1:0] ram_w32_l128_id11_1_addr,
  output [32-1:0] ram_w32_l128_id11_1_rdata,
  input [32-1:0] ram_w32_l128_id11_1_wdata,
  input ram_w32_l128_id11_1_wenable,
  input ram_w32_l128_id11_1_enable
);

  reg [32-1:0] ram_w32_l128_id11_0_rdata_out;
  assign ram_w32_l128_id11_0_rdata = ram_w32_l128_id11_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id11_1_rdata_out;
  assign ram_w32_l128_id11_1_rdata = ram_w32_l128_id11_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id11_0_enable) begin
      if(ram_w32_l128_id11_0_wenable) begin
        mem[ram_w32_l128_id11_0_addr] <= ram_w32_l128_id11_0_wdata;
        ram_w32_l128_id11_0_rdata_out <= ram_w32_l128_id11_0_wdata;
      end else begin
        ram_w32_l128_id11_0_rdata_out <= mem[ram_w32_l128_id11_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id11_1_enable) begin
      if(ram_w32_l128_id11_1_wenable) begin
        mem[ram_w32_l128_id11_1_addr] <= ram_w32_l128_id11_1_wdata;
        ram_w32_l128_id11_1_rdata_out <= ram_w32_l128_id11_1_wdata;
      end else begin
        ram_w32_l128_id11_1_rdata_out <= mem[ram_w32_l128_id11_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id12
(
  input CLK,
  input [7-1:0] ram_w32_l128_id12_0_addr,
  output [32-1:0] ram_w32_l128_id12_0_rdata,
  input [32-1:0] ram_w32_l128_id12_0_wdata,
  input ram_w32_l128_id12_0_wenable,
  input ram_w32_l128_id12_0_enable,
  input [7-1:0] ram_w32_l128_id12_1_addr,
  output [32-1:0] ram_w32_l128_id12_1_rdata,
  input [32-1:0] ram_w32_l128_id12_1_wdata,
  input ram_w32_l128_id12_1_wenable,
  input ram_w32_l128_id12_1_enable
);

  reg [32-1:0] ram_w32_l128_id12_0_rdata_out;
  assign ram_w32_l128_id12_0_rdata = ram_w32_l128_id12_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id12_1_rdata_out;
  assign ram_w32_l128_id12_1_rdata = ram_w32_l128_id12_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id12_0_enable) begin
      if(ram_w32_l128_id12_0_wenable) begin
        mem[ram_w32_l128_id12_0_addr] <= ram_w32_l128_id12_0_wdata;
        ram_w32_l128_id12_0_rdata_out <= ram_w32_l128_id12_0_wdata;
      end else begin
        ram_w32_l128_id12_0_rdata_out <= mem[ram_w32_l128_id12_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id12_1_enable) begin
      if(ram_w32_l128_id12_1_wenable) begin
        mem[ram_w32_l128_id12_1_addr] <= ram_w32_l128_id12_1_wdata;
        ram_w32_l128_id12_1_rdata_out <= ram_w32_l128_id12_1_wdata;
      end else begin
        ram_w32_l128_id12_1_rdata_out <= mem[ram_w32_l128_id12_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id13
(
  input CLK,
  input [7-1:0] ram_w32_l128_id13_0_addr,
  output [32-1:0] ram_w32_l128_id13_0_rdata,
  input [32-1:0] ram_w32_l128_id13_0_wdata,
  input ram_w32_l128_id13_0_wenable,
  input ram_w32_l128_id13_0_enable,
  input [7-1:0] ram_w32_l128_id13_1_addr,
  output [32-1:0] ram_w32_l128_id13_1_rdata,
  input [32-1:0] ram_w32_l128_id13_1_wdata,
  input ram_w32_l128_id13_1_wenable,
  input ram_w32_l128_id13_1_enable
);

  reg [32-1:0] ram_w32_l128_id13_0_rdata_out;
  assign ram_w32_l128_id13_0_rdata = ram_w32_l128_id13_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id13_1_rdata_out;
  assign ram_w32_l128_id13_1_rdata = ram_w32_l128_id13_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id13_0_enable) begin
      if(ram_w32_l128_id13_0_wenable) begin
        mem[ram_w32_l128_id13_0_addr] <= ram_w32_l128_id13_0_wdata;
        ram_w32_l128_id13_0_rdata_out <= ram_w32_l128_id13_0_wdata;
      end else begin
        ram_w32_l128_id13_0_rdata_out <= mem[ram_w32_l128_id13_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id13_1_enable) begin
      if(ram_w32_l128_id13_1_wenable) begin
        mem[ram_w32_l128_id13_1_addr] <= ram_w32_l128_id13_1_wdata;
        ram_w32_l128_id13_1_rdata_out <= ram_w32_l128_id13_1_wdata;
      end else begin
        ram_w32_l128_id13_1_rdata_out <= mem[ram_w32_l128_id13_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id14
(
  input CLK,
  input [7-1:0] ram_w32_l128_id14_0_addr,
  output [32-1:0] ram_w32_l128_id14_0_rdata,
  input [32-1:0] ram_w32_l128_id14_0_wdata,
  input ram_w32_l128_id14_0_wenable,
  input ram_w32_l128_id14_0_enable,
  input [7-1:0] ram_w32_l128_id14_1_addr,
  output [32-1:0] ram_w32_l128_id14_1_rdata,
  input [32-1:0] ram_w32_l128_id14_1_wdata,
  input ram_w32_l128_id14_1_wenable,
  input ram_w32_l128_id14_1_enable
);

  reg [32-1:0] ram_w32_l128_id14_0_rdata_out;
  assign ram_w32_l128_id14_0_rdata = ram_w32_l128_id14_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id14_1_rdata_out;
  assign ram_w32_l128_id14_1_rdata = ram_w32_l128_id14_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id14_0_enable) begin
      if(ram_w32_l128_id14_0_wenable) begin
        mem[ram_w32_l128_id14_0_addr] <= ram_w32_l128_id14_0_wdata;
        ram_w32_l128_id14_0_rdata_out <= ram_w32_l128_id14_0_wdata;
      end else begin
        ram_w32_l128_id14_0_rdata_out <= mem[ram_w32_l128_id14_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id14_1_enable) begin
      if(ram_w32_l128_id14_1_wenable) begin
        mem[ram_w32_l128_id14_1_addr] <= ram_w32_l128_id14_1_wdata;
        ram_w32_l128_id14_1_rdata_out <= ram_w32_l128_id14_1_wdata;
      end else begin
        ram_w32_l128_id14_1_rdata_out <= mem[ram_w32_l128_id14_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id15
(
  input CLK,
  input [7-1:0] ram_w32_l128_id15_0_addr,
  output [32-1:0] ram_w32_l128_id15_0_rdata,
  input [32-1:0] ram_w32_l128_id15_0_wdata,
  input ram_w32_l128_id15_0_wenable,
  input ram_w32_l128_id15_0_enable,
  input [7-1:0] ram_w32_l128_id15_1_addr,
  output [32-1:0] ram_w32_l128_id15_1_rdata,
  input [32-1:0] ram_w32_l128_id15_1_wdata,
  input ram_w32_l128_id15_1_wenable,
  input ram_w32_l128_id15_1_enable
);

  reg [32-1:0] ram_w32_l128_id15_0_rdata_out;
  assign ram_w32_l128_id15_0_rdata = ram_w32_l128_id15_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id15_1_rdata_out;
  assign ram_w32_l128_id15_1_rdata = ram_w32_l128_id15_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id15_0_enable) begin
      if(ram_w32_l128_id15_0_wenable) begin
        mem[ram_w32_l128_id15_0_addr] <= ram_w32_l128_id15_0_wdata;
        ram_w32_l128_id15_0_rdata_out <= ram_w32_l128_id15_0_wdata;
      end else begin
        ram_w32_l128_id15_0_rdata_out <= mem[ram_w32_l128_id15_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id15_1_enable) begin
      if(ram_w32_l128_id15_1_wenable) begin
        mem[ram_w32_l128_id15_1_addr] <= ram_w32_l128_id15_1_wdata;
        ram_w32_l128_id15_1_rdata_out <= ram_w32_l128_id15_1_wdata;
      end else begin
        ram_w32_l128_id15_1_rdata_out <= mem[ram_w32_l128_id15_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id16
(
  input CLK,
  input [7-1:0] ram_w32_l128_id16_0_addr,
  output [32-1:0] ram_w32_l128_id16_0_rdata,
  input [32-1:0] ram_w32_l128_id16_0_wdata,
  input ram_w32_l128_id16_0_wenable,
  input ram_w32_l128_id16_0_enable,
  input [7-1:0] ram_w32_l128_id16_1_addr,
  output [32-1:0] ram_w32_l128_id16_1_rdata,
  input [32-1:0] ram_w32_l128_id16_1_wdata,
  input ram_w32_l128_id16_1_wenable,
  input ram_w32_l128_id16_1_enable
);

  reg [32-1:0] ram_w32_l128_id16_0_rdata_out;
  assign ram_w32_l128_id16_0_rdata = ram_w32_l128_id16_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id16_1_rdata_out;
  assign ram_w32_l128_id16_1_rdata = ram_w32_l128_id16_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id16_0_enable) begin
      if(ram_w32_l128_id16_0_wenable) begin
        mem[ram_w32_l128_id16_0_addr] <= ram_w32_l128_id16_0_wdata;
        ram_w32_l128_id16_0_rdata_out <= ram_w32_l128_id16_0_wdata;
      end else begin
        ram_w32_l128_id16_0_rdata_out <= mem[ram_w32_l128_id16_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id16_1_enable) begin
      if(ram_w32_l128_id16_1_wenable) begin
        mem[ram_w32_l128_id16_1_addr] <= ram_w32_l128_id16_1_wdata;
        ram_w32_l128_id16_1_rdata_out <= ram_w32_l128_id16_1_wdata;
      end else begin
        ram_w32_l128_id16_1_rdata_out <= mem[ram_w32_l128_id16_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id17
(
  input CLK,
  input [7-1:0] ram_w32_l128_id17_0_addr,
  output [32-1:0] ram_w32_l128_id17_0_rdata,
  input [32-1:0] ram_w32_l128_id17_0_wdata,
  input ram_w32_l128_id17_0_wenable,
  input ram_w32_l128_id17_0_enable,
  input [7-1:0] ram_w32_l128_id17_1_addr,
  output [32-1:0] ram_w32_l128_id17_1_rdata,
  input [32-1:0] ram_w32_l128_id17_1_wdata,
  input ram_w32_l128_id17_1_wenable,
  input ram_w32_l128_id17_1_enable
);

  reg [32-1:0] ram_w32_l128_id17_0_rdata_out;
  assign ram_w32_l128_id17_0_rdata = ram_w32_l128_id17_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id17_1_rdata_out;
  assign ram_w32_l128_id17_1_rdata = ram_w32_l128_id17_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id17_0_enable) begin
      if(ram_w32_l128_id17_0_wenable) begin
        mem[ram_w32_l128_id17_0_addr] <= ram_w32_l128_id17_0_wdata;
        ram_w32_l128_id17_0_rdata_out <= ram_w32_l128_id17_0_wdata;
      end else begin
        ram_w32_l128_id17_0_rdata_out <= mem[ram_w32_l128_id17_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id17_1_enable) begin
      if(ram_w32_l128_id17_1_wenable) begin
        mem[ram_w32_l128_id17_1_addr] <= ram_w32_l128_id17_1_wdata;
        ram_w32_l128_id17_1_rdata_out <= ram_w32_l128_id17_1_wdata;
      end else begin
        ram_w32_l128_id17_1_rdata_out <= mem[ram_w32_l128_id17_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l128_id18
(
  input CLK,
  input [7-1:0] ram_w32_l128_id18_0_addr,
  output [32-1:0] ram_w32_l128_id18_0_rdata,
  input [32-1:0] ram_w32_l128_id18_0_wdata,
  input ram_w32_l128_id18_0_wenable,
  input ram_w32_l128_id18_0_enable,
  input [7-1:0] ram_w32_l128_id18_1_addr,
  output [32-1:0] ram_w32_l128_id18_1_rdata,
  input [32-1:0] ram_w32_l128_id18_1_wdata,
  input ram_w32_l128_id18_1_wenable,
  input ram_w32_l128_id18_1_enable
);

  reg [32-1:0] ram_w32_l128_id18_0_rdata_out;
  assign ram_w32_l128_id18_0_rdata = ram_w32_l128_id18_0_rdata_out;
  reg [32-1:0] ram_w32_l128_id18_1_rdata_out;
  assign ram_w32_l128_id18_1_rdata = ram_w32_l128_id18_1_rdata_out;
  reg [32-1:0] mem [0:128-1];

  always @(posedge CLK) begin
    if(ram_w32_l128_id18_0_enable) begin
      if(ram_w32_l128_id18_0_wenable) begin
        mem[ram_w32_l128_id18_0_addr] <= ram_w32_l128_id18_0_wdata;
        ram_w32_l128_id18_0_rdata_out <= ram_w32_l128_id18_0_wdata;
      end else begin
        ram_w32_l128_id18_0_rdata_out <= mem[ram_w32_l128_id18_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l128_id18_1_enable) begin
      if(ram_w32_l128_id18_1_wenable) begin
        mem[ram_w32_l128_id18_1_addr] <= ram_w32_l128_id18_1_wdata;
        ram_w32_l128_id18_1_rdata_out <= ram_w32_l128_id18_1_wdata;
      end else begin
        ram_w32_l128_id18_1_rdata_out <= mem[ram_w32_l128_id18_1_addr];
      end
    end 
  end


endmodule



module madd_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_0
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_1
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_2
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_2
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_2
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_3
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_3
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_3
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_4
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_4
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_4
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_5
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_5
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_5
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_6
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_6
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_6
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_7
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_7
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_7
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_8
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_8
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_8
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  output [64-1:0] c
);


  multiplier_core_0
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  output [64-1:0] c
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  wire signed [64-1:0] _mul;
  reg signed [64-1:0] _pipe_mul0;
  reg signed [64-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule



module multiplier_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [7-1:0] b,
  output [39-1:0] c
);


  multiplier_core_1
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [7-1:0] b,
  output [39-1:0] c
);

  reg signed [32-1:0] _a;
  reg signed [7-1:0] _b;
  wire signed [39-1:0] _mul;
  reg signed [39-1:0] _pipe_mul0;
  assign _mul = _a * _b;
  assign c = _pipe_mul0;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
    end 
  end


endmodule



module _lut_LUT_ROM_857
(
  input CLK,
  input [8-1:0] addr,
  input enable,
  output reg [32-1:0] val
);


  always @(posedge CLK) begin
    if(enable) begin
      case(addr)
        0: begin
          val <= 0;
        end
        1: begin
          val <= -49746405;
        end
        2: begin
          val <= -98340436;
        end
        3: begin
          val <= -145808787;
        end
        4: begin
          val <= -192177536;
        end
        5: begin
          val <= -237472153;
        end
        6: begin
          val <= -281717522;
        end
        7: begin
          val <= -324937947;
        end
        8: begin
          val <= -367157173;
        end
        9: begin
          val <= -408398391;
        end
        10: begin
          val <= -448684258;
        end
        11: begin
          val <= -488036903;
        end
        12: begin
          val <= -526477946;
        end
        13: begin
          val <= -564028503;
        end
        14: begin
          val <= -600709201;
        end
        15: begin
          val <= -636540193;
        end
        16: begin
          val <= -671541160;
        end
        17: begin
          val <= -705731331;
        end
        18: begin
          val <= -739129488;
        end
        19: begin
          val <= -771753977;
        end
        20: begin
          val <= -803622720;
        end
        21: begin
          val <= -834753225;
        end
        22: begin
          val <= -865162593;
        end
        23: begin
          val <= -894867528;
        end
        24: begin
          val <= -923884349;
        end
        25: begin
          val <= -952228996;
        end
        26: begin
          val <= -979917040;
        end
        27: begin
          val <= -1006963692;
        end
        28: begin
          val <= -1033383808;
        end
        29: begin
          val <= -1059191903;
        end
        30: begin
          val <= -1084402154;
        end
        31: begin
          val <= -1109028410;
        end
        32: begin
          val <= -1133084200;
        end
        33: begin
          val <= -1156582738;
        end
        34: begin
          val <= -1179536933;
        end
        35: begin
          val <= -1201959394;
        end
        36: begin
          val <= -1223862440;
        end
        37: begin
          val <= -1245258102;
        end
        38: begin
          val <= -1266158135;
        end
        39: begin
          val <= -1286574018;
        end
        40: begin
          val <= -1306516968;
        end
        41: begin
          val <= -1325997940;
        end
        42: begin
          val <= -1345027636;
        end
        43: begin
          val <= -1363616510;
        end
        44: begin
          val <= -1381774773;
        end
        45: begin
          val <= -1399512400;
        end
        46: begin
          val <= -1416839135;
        end
        47: begin
          val <= -1433764497;
        end
        48: begin
          val <= -1450297783;
        end
        49: begin
          val <= -1466448076;
        end
        50: begin
          val <= -1482224248;
        end
        51: begin
          val <= -1497634966;
        end
        52: begin
          val <= -1512688694;
        end
        53: begin
          val <= -1527393703;
        end
        54: begin
          val <= -1541758072;
        end
        55: begin
          val <= -1555789689;
        end
        56: begin
          val <= -1569496265;
        end
        57: begin
          val <= -1582885328;
        end
        58: begin
          val <= -1595964234;
        end
        59: begin
          val <= -1608740168;
        end
        60: begin
          val <= -1621220147;
        end
        61: begin
          val <= -1633411028;
        end
        62: begin
          val <= -1645319507;
        end
        63: begin
          val <= -1656952127;
        end
        64: begin
          val <= -1668315278;
        end
        65: begin
          val <= -1679415201;
        end
        66: begin
          val <= -1690257995;
        end
        67: begin
          val <= -1700849616;
        end
        68: begin
          val <= -1711195882;
        end
        69: begin
          val <= -1721302477;
        end
        70: begin
          val <= -1731174953;
        end
        71: begin
          val <= -1740818734;
        end
        72: begin
          val <= -1750239117;
        end
        73: begin
          val <= -1759441276;
        end
        74: begin
          val <= -1768430268;
        end
        75: begin
          val <= -1777211030;
        end
        76: begin
          val <= -1785788386;
        end
        77: begin
          val <= -1794167048;
        end
        78: begin
          val <= -1802351618;
        end
        79: begin
          val <= -1810346593;
        end
        80: begin
          val <= -1818156364;
        end
        81: begin
          val <= -1825785223;
        end
        82: begin
          val <= -1833237359;
        end
        83: begin
          val <= -1840516866;
        end
        84: begin
          val <= -1847627744;
        end
        85: begin
          val <= -1854573898;
        end
        86: begin
          val <= -1861359146;
        end
        87: begin
          val <= -1867987212;
        end
        88: begin
          val <= -1874461740;
        end
        89: begin
          val <= -1880786286;
        end
        90: begin
          val <= -1886964324;
        end
        91: begin
          val <= -1892999248;
        end
        92: begin
          val <= -1898894372;
        end
        93: begin
          val <= -1904652937;
        end
        94: begin
          val <= -1910278104;
        end
        95: begin
          val <= -1915772965;
        end
        96: begin
          val <= -1921140537;
        end
        97: begin
          val <= -1926383769;
        end
        98: begin
          val <= -1931505542;
        end
        99: begin
          val <= -1936508670;
        end
        100: begin
          val <= -1941395900;
        end
        101: begin
          val <= -1946169918;
        end
        102: begin
          val <= -1950833345;
        end
        103: begin
          val <= -1955388744;
        end
        104: begin
          val <= -1959838618;
        end
        105: begin
          val <= -1964185411;
        end
        106: begin
          val <= -1968431510;
        end
        107: begin
          val <= -1972579248;
        end
        108: begin
          val <= -1976630904;
        end
        109: begin
          val <= -1980588704;
        end
        110: begin
          val <= -1984454821;
        end
        111: begin
          val <= -1988231379;
        end
        112: begin
          val <= -1991920454;
        end
        113: begin
          val <= -1995524072;
        end
        114: begin
          val <= -1999044212;
        end
        115: begin
          val <= -2002482807;
        end
        116: begin
          val <= -2005841748;
        end
        117: begin
          val <= -2009122879;
        end
        118: begin
          val <= -2012328003;
        end
        119: begin
          val <= -2015458880;
        end
        120: begin
          val <= -2018517231;
        end
        121: begin
          val <= -2021504735;
        end
        122: begin
          val <= -2024423033;
        end
        123: begin
          val <= -2027273729;
        end
        124: begin
          val <= -2030058389;
        end
        125: begin
          val <= -2032778542;
        end
        126: begin
          val <= -2035435683;
        end
        127: begin
          val <= -2038031271;
        end
        128: begin
          val <= -2040566733;
        end
        129: begin
          val <= -2043043460;
        end
        130: begin
          val <= -2045462815;
        end
        131: begin
          val <= -2047826125;
        end
        132: begin
          val <= -2050134689;
        end
        133: begin
          val <= -2052389775;
        end
        134: begin
          val <= -2054592622;
        end
        135: begin
          val <= -2056744441;
        end
        136: begin
          val <= -2058846412;
        end
        137: begin
          val <= -2060899691;
        end
        138: begin
          val <= -2062905407;
        end
        139: begin
          val <= -2064864659;
        end
        140: begin
          val <= -2066778526;
        end
        141: begin
          val <= -2068648058;
        end
        142: begin
          val <= -2070474283;
        end
        143: begin
          val <= -2072258203;
        end
        144: begin
          val <= -2074000798;
        end
        145: begin
          val <= -2075703027;
        end
        146: begin
          val <= -2077365823;
        end
        147: begin
          val <= -2078990101;
        end
        148: begin
          val <= -2080576752;
        end
        149: begin
          val <= -2082126649;
        end
        150: begin
          val <= -2083640642;
        end
        151: begin
          val <= -2085119564;
        end
        152: begin
          val <= -2086564226;
        end
        153: begin
          val <= -2087975423;
        end
        154: begin
          val <= -2089353929;
        end
        155: begin
          val <= -2090700503;
        end
        156: begin
          val <= -2092015883;
        end
        157: begin
          val <= -2093300792;
        end
        158: begin
          val <= -2094555937;
        end
        159: begin
          val <= -2095782006;
        end
        160: begin
          val <= -2096979673;
        end
        161: begin
          val <= -2098149597;
        end
        162: begin
          val <= -2099292419;
        end
        163: begin
          val <= -2100408767;
        end
        164: begin
          val <= -2101499256;
        end
        165: begin
          val <= -2102564483;
        end
        166: begin
          val <= -2103605034;
        end
        167: begin
          val <= -2104621481;
        end
        168: begin
          val <= -2105614382;
        end
        169: begin
          val <= -2106584283;
        end
        170: begin
          val <= -2107531716;
        end
        171: begin
          val <= -2108457201;
        end
        172: begin
          val <= -2109361248;
        end
        173: begin
          val <= -2110244352;
        end
        174: begin
          val <= -2111107000;
        end
        175: begin
          val <= -2111949664;
        end
        176: begin
          val <= -2112772808;
        end
        177: begin
          val <= -2113576883;
        end
        178: begin
          val <= -2114362333;
        end
        179: begin
          val <= -2115129587;
        end
        180: begin
          val <= -2115879068;
        end
        181: begin
          val <= -2116611188;
        end
        182: begin
          val <= -2117326347;
        end
        183: begin
          val <= -2118024940;
        end
        184: begin
          val <= -2118707351;
        end
        185: begin
          val <= -2119373953;
        end
        186: begin
          val <= -2120025113;
        end
        187: begin
          val <= -2120661190;
        end
        188: begin
          val <= -2121282531;
        end
        189: begin
          val <= -2121889479;
        end
        190: begin
          val <= -2122482368;
        end
        191: begin
          val <= -2123061522;
        end
        192: begin
          val <= -2123627260;
        end
        193: begin
          val <= -2124179892;
        end
        194: begin
          val <= -2124719723;
        end
        195: begin
          val <= -2125247049;
        end
        196: begin
          val <= -2125762159;
        end
        197: begin
          val <= -2126265337;
        end
        198: begin
          val <= -2126756859;
        end
        199: begin
          val <= -2127236994;
        end
        200: begin
          val <= -2127706007;
        end
        201: begin
          val <= -2128164156;
        end
        202: begin
          val <= -2128611691;
        end
        203: begin
          val <= -2129048860;
        end
        204: begin
          val <= -2129475901;
        end
        205: begin
          val <= -2129893050;
        end
        206: begin
          val <= -2130300536;
        end
        207: begin
          val <= -2130698582;
        end
        208: begin
          val <= -2131087408;
        end
        209: begin
          val <= -2131467227;
        end
        210: begin
          val <= -2131838247;
        end
        211: begin
          val <= -2132200672;
        end
        212: begin
          val <= -2132554702;
        end
        213: begin
          val <= -2132900530;
        end
        214: begin
          val <= -2133238348;
        end
        215: begin
          val <= -2133568340;
        end
        216: begin
          val <= -2133890688;
        end
        217: begin
          val <= -2134205568;
        end
        218: begin
          val <= -2134513155;
        end
        219: begin
          val <= -2134813616;
        end
        220: begin
          val <= -2135107117;
        end
        221: begin
          val <= -2135393819;
        end
        222: begin
          val <= -2135673879;
        end
        223: begin
          val <= -2135947452;
        end
        224: begin
          val <= -2136214688;
        end
        225: begin
          val <= -2136475733;
        end
        226: begin
          val <= -2136730731;
        end
        227: begin
          val <= -2136979822;
        end
        228: begin
          val <= -2137223143;
        end
        229: begin
          val <= -2137460828;
        end
        230: begin
          val <= -2137693006;
        end
        231: begin
          val <= -2137919806;
        end
        232: begin
          val <= -2138141352;
        end
        233: begin
          val <= -2138357766;
        end
        234: begin
          val <= -2138569167;
        end
        235: begin
          val <= -2138775671;
        end
        236: begin
          val <= -2138977391;
        end
        237: begin
          val <= -2139174438;
        end
        238: begin
          val <= -2139366921;
        end
        239: begin
          val <= -2139554944;
        end
        240: begin
          val <= -2139738613;
        end
        241: begin
          val <= -2139918026;
        end
        242: begin
          val <= -2140093284;
        end
        243: begin
          val <= -2140264481;
        end
        244: begin
          val <= -2140431713;
        end
        245: begin
          val <= -2140595071;
        end
        246: begin
          val <= -2140754645;
        end
        247: begin
          val <= -2140910522;
        end
        248: begin
          val <= -2141062788;
        end
        249: begin
          val <= -2141211527;
        end
        250: begin
          val <= -2141356821;
        end
        251: begin
          val <= -2141498749;
        end
        252: begin
          val <= -2141637389;
        end
        253: begin
          val <= -2141772817;
        end
        254: begin
          val <= -2141905108;
        end
        255: begin
          val <= -2142034335;
        end
      endcase
    end 
  end


endmodule

